��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��g��C�$	��&�1�noX�j y�{���(�����:]�2 ��lY.�~H�+�"�yfA�H5RDY�8�R�*z��r��a�TG f;+�:��V���3/O�u�0��*�N������-���a������3{�$\x �_�T��Qo6(��t�s�����{�p�� O	��[�zɜZ�v6]�b׼�e�*��5�U)�)��y�/\�xpR幎n���J�V��V&��]W�S��V�w��y\���D]Ȋn�(D��,�B7p%�/�AsI�X����Uh$ip�C�[E2��Ӟ�&.��lu���.��&ùU>���r�
��kO]S>y�(�g���t0�l�����ʭ�Vs���2��`M��>�H�y�is��(i<�������=����C��{��	M�{�x�]�l9�nfǿ��E���yDs�9��o�!��Q�8���aY��AKv���%Gj��so�#�[EEd�L�����j+{\���{�[2`��54�f��3�C��/S���7�	���M�C���f�G��*���0ؾ� S��6p]�@���4BBjg���o�3���h��0�Gۮ��:����b�)�/9I�D�g��`c�@ez{��,�!d���=�Ka�7=i���^t��U����"��gP��EE3�,De�5Shd��k����_������B����=x��tG��J���]�%�`�<�vtUHܸ�W���t.'�����5G�D;S��V�r
V,�aBZ���d��lX
���Ұ8�L��}�?��S3��Ts����x\�O�V�w��c�?<��1�44e������Lǚe&��Ŷw]F��
x
�9`��۶zQBX�A�
�	��z���&}���$|�.���O���(�ۤ9��e7`��`Qr�&�+
(P%g��0��� P��gY�:������͌}�%�L�o����붞�`B��f���5�:%e,�@S�7����g>���~K~5����
?�fLzrGJ�a�"���9;D��wRU���;��$M�A/B�K@ʌ�<*�a�5�yMi���4p�n1��������am���`�m���E\�R�r���F��ԑ�@J�J)վF���q���X>:��	Q
 e&&.5�o�^<�l��	��B��C�+$h)u��t(��7L��ʆ\��	��L�f^H�ԍoە�焙��>Ns�Yl8��Atﲲs�����k�r#U�&W�G���X��(���edY;��Ç����a�fL�Paί����?��p2D�k~1���,4��v]{��s�Z�b�<�̣�Ġ��:�������X:x�����X�&%TC�Ҽ���}��6��A.sҬN���v�B���fg���S�-�4������Ĩ1��^41��X���fO��^�{����!�\+�a��(�I]	�Vp�cJ�uT*W��;=���9�GheU_���R�,W���8�ZR��
��x�3C�o�G��0"Bom�C9M����ĉ�d���Yc�Lr��"����,G��0M�U��k�fZ-��й�M��ٻ�j$����L������j@�N����5�h1������@߁���J@HbIU��ي���:�,�o|��zI�ak��7&��>�� �+MXֲA�
�<�z��z��K�U�=���.v��Z({�3������o�od�3i�Ї�[>y'd?�k9I/i�#>~�`�T��<�d\�)���F��c�5�ǻ;"Ɔ����&�����A�uR�Qݮ�Ï���&�No!,����������>�e��1}I�Q�w~Q�v	���Qة��F_R�魮�M�3�>�X2�W�B�@*g��`!���E��e)��n)/�3�"�(|�F���`V��
��N�^B9�a���'�����w��C�z8ݰ�Ü4����e����¡�aJ��#��N1��t$>4ﯨ��MwB��H��X�i�B��Ghe0/b�3N�X,����f�}]�����f�G��|�=ݠ��2=����V$@_�K����=>76�g�[OXؓ*U�`qs��.��K�c�S�nu�)d�x��<��p����I����<<��ǔ�5��$?�r�o:1����+�o�'��5���!(PceW��)O`��8IE�󽙕A����]4�A�'�c�'}ݿ���J�-�<��R젘�1���J����	J��3�` qJk�. ���%!l������7���8"�ƚ6ԣBҴ�T�*��q�&R �Ye��V[����+���ǜpN��9	��}�p33r���P��ҷ�v
���[ĉ6LM���_itj����T�|k������\��8�XQ4�bgV���V���i%!��sݗ�k� i#Ώ���H�L5U�y�Ext��ٴ� �qo���mK�1�	m��k|��z;b�EQl���wfz�#��7wKD�߻�x&��բW�ԤQSv�Ԋ|���s����}r�_\��`���5�c�����>jmGXI�b�g5�
3�*��F�qۼ��lP3:q�����r�����j�j��{aj���20c�V
HXo�r��_������*�j3��_�f<��<�?�Ez"�D��=���� ޱ$G���L@����Oi�g�"����Te qE��kWz�#$��`:����DM]N8e1�PY����R�6'��\V��/����]��6�c��K%1��B���#:�m�Wѭ�5�7�{W�s`$����h��uX��!���a������k���@��Z�L�״���(���J�W^�M�x��y���v-9��.�AY�hixN��t�Zt�d�}oT��.8\ ?�{3�[F��℩T;�G#��_8�%�����o����
��2�k��^�̳������P�n����T�P���Fde2QF����Uiʆ�,���)���pi�|�]�}fm1-�l�~)��n�}�+���	���k�;t�T�����^�gM��Nm���9W�|�PC�g\T�B/�a�D̰�l ��
��l)â�g�j�́��6�U�!�Y+lsVEO C8)�H�5�?�A'+kMF���,G��t��bQ� �,@�������1q�t��PR�^�����D`��H3��h���.[��x�D�NY�oW�T�#6�N����ނ���_��"?�kz�q�(�qSvVŃ죢=��CƐ�4�]�{�W��,�Pb:ۆ_�O!�`ѷ�2���Ѭ�`ꅸ�������׹�S�d�%�/���]r��<��Ӥ�z�Rb�mh�ȝ��}jFP("^X���<~�O�0O=��b�orO����[R]��q`4~�:��� zϪV(z��9_E�V����\H�Ī�oj��(e�����l�����P�b�yŎ5�(
��u�_-?�M����B%aQ�:_鑕�ɵJ��x���Z�c�ؾ��	�?�w�����.��4B�)9��#��G���4�����<["�o�� oH{��]f�rY�FR�FF#t0%��~v4���E�ٔ[�vv�w� ����lT�1�p���+��p�
:ßU)��CHj|��h'��j��?L>N��T��U�Կ���KK��6=h`��u�����{^6��p	qR5���ь�6�A�i-���nBD�lkN=��_Na_>�$g��X�<^w9������+�z���m�� ��`������=��vi0�KB>�J�Y@-�i���Ŀ1��7ehetz4�%n��ƽ���ݟ?���ew�Sו��d`V�+�-~��c�j��KM����Oi��(����=�gо�����
�s���1������Ų�(�j�3��Ǟ)�Q<�$X�.D�9�*�9[�Qf��gF�9A+�Օ�'�#���/=棭�{"�Y�ԠT���JtU�:�V� �
_���b+rz���y'.��$@�z)Пf�l�3�v)Dc��)oq�(s&b�nΜ��G�o�(�<�A��{5ZnZ&x�_������P����'T ����3�Ww�L!=� m8e@.�s�.�=kAզtRP��y�e�%Q�*>r��ya�P�ENl0���V*��T�ǡ;`[�f�L�|��ռ�����J��=o�É[���%�g��|0a@�`�7m��$�[%��Q��]ߋ�E���( ���l����O2scC��oR��N��W�'�=^0�;�=�o�a:��+ЬB���=^�τ��6�˄h�K��;� ���`<�T��	�}��N� �z�E��DsڡN<G���F���D��������@�K�#q�!�*�mn�����y�jR�H�����̶^F�Z[�:AW����3bBsbj�[�e���c	�aD�@��:��՝#3����Ra��8�צ�K���R�D��X�qk�(�t��@�K�T#��P!M0�(��5m����E���e��Gp�t�����\:s�{�m��H�t`�i�0H���$2�[�pR���NA���V~��vO��u���ژD��2��T1�w�!r��/����H���8������킙�3zz���4�1D��<��u��Xg�@�(�$\yȘ4�|BEtX���'ֻ�T�p��[�|���I8�5@H��0��(��ܐ�R�L�$�df�V���h:���=Rs�P��b��><	ʴ,���S�YU�z�����YT鿏�N*�N\F��~N���~;ya*[���c���Zh��J��s}���4Eć���9�����#�@���[x�����$ӄs�l<�<�pd�*}֝@��=zlF R�����n�I�K�,�B{��O�1$�}��p3*tޑ r�t�w���_�V�=�����M�=Q�4;�x�L��E{c��?�hq�1��~��������#�TBobGR�w��"ą�ee@��S kx(�G���HX�~�	\�T�7l��C��H����{zh��A����Η50�=��K|f�H�2�|l�P�9 C�z���\�s"��]d'4as�b�G��j�m���>"i�Q��\CXS"��}Í(��/=ە*�������~X&������6��4e�Uq�6��N����N��V��7s�!>op 2�z�n��6mm�GYE��?��٬�I�X���_��Ut�6�A�eR��`���QJSHb�b,������2K�x���H���Ka|�}]��К?��蓃���Fd/I[8R��R�s��y����E-��
K�����{��b���o��C�>v�8�,��\�����6s�`<�7����g,�n	�j�A�K;�]��tK�|pglj|@y�L��Y+�����/��H�v4Bǹq8?�>�B�S*�%ۺi��K�N���M4��%�?HZ]���%k������O�Nmjo�`���m3���d���x�6G��C���c(�w4���\�ԕIF��z�%�:��e�YV�gg�tt�����f��ؾ
��xߴ)��l��{}i���d��G�,��B��!Pt@�u���(��]`.�������Ix'#b����_�X�P� ���:����5�93�qJ��%3â2QA�Pn!��uĞ!C���UCi"�~#i�qR0s�U��`����PQ���L�E
����4��KD�~�u�g�c���]X��fQ�������[f��	(O�%SϏ?�����6:�����ޗ$X�%�{Ro��1��p�<*.�-Ӽ����[<��M���9'nrj�tK��8�+�C��(�BV˒X��d�
l�	@�3�����.�
��py����!�� ��
D���D�*��=���1��?Y�+���o�r�
�2MJ�x��4K��z�Ci��gw��Y��X�&�^������n7��@~<���E��5��d�uWcw�Y�9讬m[:��1����3�_�bU�ږ���DQ�-��-/��K7�(D %��3=�d�^8���jW��+��*U�K����w���\��/�Fct86�Y<�\� ����Ū>ך�\�@*��}#f��Y�V/"��v,�F^������C�����P�V��lkr1,Y�qbTy��# �2�g���gsi�E�GV�(��& ���I���&_tx�K�\��U���kz�Ƨ���K�9_��%�T�?���&�w��/�e��[�>F�L�$`��%��Q��}�;���&�0��江��1>X��_�T��`�TJ���Ea2�]YjX��s3ʏ��N��f2@����1�(�Ւ
A�z2�ʰ���#�]��[��o-G�u�=E�	��]�I���qN���W�Z|�E�"4�����N�v�_P��B!�.�6����
�}���+�`��F�P]x�IG�h_*�>�)ڠ���[\�?H�� ��}$.4/.�z�>Wk�Ĵ�y�r�[W'����jn��;�i�-Pi�d��8`�m�1�z�ݹ ����aTn>�Yl�	^u�1:���%E�J&��$�@|��Ӓ������'��h ߓ�4)I9w�8;��"�l!��k	����6�KB�vPmp^|�\ǚP��[�!d���aZ6푉��)͵��bl�Vx�:�gy ~�U0b�4~Z_X�q"Z��KTߪ��z�~��A�Q�P�9 �kJ�77'�C�1���t�(W�>��O��.�Fbs�nj\���#���#{W�0��R��
E����M�TZRa7R�}�p�����f X7 ��]����KhJa[�Z*�/�HUP �(ו��ҫJ>�u�ח��=����N�3h�x��Ś�T@Ux�@v`�%�]!cT.ͺ>bB��70 M�@��53�4SqP�,{�_�0� ����X&F�~Ců���YH���%8�%ܵr.���&�c���3�
K׍������ty�Q�t��Zw 0㈋�=_+n1�@n���7R���gPuptV�z�����_)��E��P����Er�ì��W�j�A�7�v��~!�� HgM���U�\�[?�{���6V�[3�ᢐlf7�/��4���N b:�'��w棎=�B��Ԓh�	����%QL���!�&і���@���VC4ٗ���?���,�) 4�22�V�1�Z<��E@^�p�v*�D�]�g�
96���eMw��J���Q�sJ�s�Н)����|�4hf�dG�>�ަ��WS��bW�g������ρ��wB���X��Ҁey{�8\-����`�:)$ :�!x�Ճ��y�Mz*j��Q�A�6�1om�޿qłw�� �D�f(v�po�<��ZZuȏ�TV�����w�J�{;u�\����Oq�`�`�lOpW �Z}�N�ɪ���3
&�~�>1�nt�~�~���7���F�Д��-3B5 ���ꫧ_� ��T0zfN@����e!�>.�Q���/��at�t`J�.!�c����}\V���֐,�G9�!BQ��E�%��hc7_�Y+ņ�aʵj`<���ಣ�I�z�6�b3��b�51��z�B��!�6������9���*/�+v,���u%����W�t�Hs�l�jW*�Ƨ�H[��b�1���֐V�@�Q�� '�ϤK7+������#0�����46!ű*�M,w�ĵۘ�1Q������[��
�w��FY๩��XK,`xņ>P���m_��<�ß3��y�\���S>�60�^���r;��r�<�1�Z�y��Ry���h��Ɩ�Ü��E}���b|v�\x�XO�NO�,U���r�n���Ƶ��������){�^4�]=�[>AK����M�v������>WO�t�ꩿ=�um�h>�ʩ�s*�@}����*ٰ9M�r�~���A}Y��D�.��|,�d_UPN5��X�� \���M��͘FP=5�AG� ���iN��Њ��x�Z�6��%𜈺[�Ⱥ��/c��z����"�M +�ܥ���o*{�+��Ǯ-�����=6?��U{�̅�4�2)"���� �@Y��9ST;�C�j�(�o�j���Uo����(o}�p���]��&=r;��s4{����2��x1/������a�"� (�	�%������1?�聑y?$����o.D��� E��ծ?P�r�'�vNVH��9���Η�#��Jތ4��p�.�;*c1��٨����W�k�nq�zx�|q~�Ž�B��M�B���ޤԉL�^���QN����iҹwL!R$��'߅�8Lc����6w�|�+����,y�)Z@�������L�c��|�������s���^w>a8��K��ݹψ5섏>y+�(�ir���Q��5�B�IRL��Q��`}�n�ʤ�:B:�M�nm%�|P-�N��m�T���n��\*s�(��ʣI�9ʞ
���kzI	7�ѯvo%����|�o��k2}?��x���5�8�i=UC�s2���r��Jce��#x�'<��b1w����.��a����s���㍏��O���l�PY?��EA��j���5��YJۮ"
�@Q��ҫ�q���_%#6�x�9�=Zz6����Lq�-vT��Q�߇u��_U�}3�B�9N_/���7n���Ɩ��!=�,�1����1U��k���)����0�!x�� ?�3ӳ�᝾�=��Ӱ�����(!#l"�uQ�5��u�!<����q��p�}�m$�r�"�F�gz��prH؈B?���;��\�|["�|��yF�����n��E�ۏ�i"��r�TQza�=^�j������-x�.8�����uf��:F6k~ȑ�q�C��]7X!)	df3g)�d>�x5�S�>�:��/6�~���[��b*�Qw��T�q]3S��iA'&���$ �+N����˂�K�$�?�I�/4螧��"LĴY��Ag�A6xx�X^�UB�zzI�GR��<FZq�Qo��=�h!@��Ơw�i)C@�n�=�:��omN5��/���$%C��o�D��|�l��J���B�c3
���2�ղR�<?�7�p�� �InR-e#t	����~Iɽ+{x�`m�kDo��`�FS(�pqr�iI�a_~�vĉ��=�>�n �h��{7~
)e�q�OX�S4�U����_	���R:QD&��pK	�௽���JP=uu��ٳ�b:J���r�����-���t��0ŭ5@��٠�@��Bu6���f2��$���}c0rE&'�����j����Y/_�q̃͡��8����S��$��*���İ�\HO�1���u�t�<3ls.ε�c�O��W�SK~^����e���0���ї>�i�����C/qT�y
��C4>���j��2"�,�LN��0P��q] �S������)Y����Ɵ��?�9*�?oI�:�*Q��ZUg�:������U����d~C�Ts�|��bY�$W
� ��}�Ӈ�i�w�N�΁��D^@n��{Z�b�34~���+r�V�z7C���36��B�yb��d,sI�1�"iq�3��m�������B�j��7H2�G�~�*�v�Nvp����M�CpbAPT1�ӊc�A�?>s.��i���C�j/MY�J��A���D��E+�D�̗*pz<�dU<�*��0��M�Yp'��Mia������,bY{U)�+�Gݾ�d�I���5�w&A����ؘ=��!�M��JU6�	��E��I�{d��9C�=�W�JkH/t7��ʋ;c�!�JB�y=퇑Am�����7��r{�5�$��Auoɣ`��*gg�<Px?��-4o��C�y��s�������d���>AA���4��D���~V|�6/�D�y�n�B���H�=Vwa�����+��`f�_�����f�O��.���`__E��g�W�ě�@�C�ϙ������0��퓤�%M�½TI�¼�����k�G39��Ur�Z@�C�X
��a��U�,M�����ђb���Bز�B$s��x�z3�t5��UZ�+� `Y����S�f����ĵ&E����ݮH����ad�f-¨�ݓ�$�/�I����� T�YEG��k �L3�(�IB��Z����E骹.��U��K[{�ʵ� �E�� �@Q8�+e��WUA������lem��45� ��l➮^%c;����A��t	8��yL�v���.
$ꢗ'צ
Ѯ�c)�7!x�7�`<�:�z�ݵ�'CT�WԦ��z5�R�]��z=����_h�)_�J�3�+G��u_ k�܊/8= si���`���CV#���殻djR�v:�PElڔ����g�����.O�L⍻ҽ7���z��%n�=���/�Ѷ��xՀp��ϕ�����f�̯�9;m���묵���u�1(£l�]σ~����a�p�d�J���h�>�F�H|l!{T����_V��k�^^�A�rFp���+�_D�W�$�K��/
'IȜI���L����˽���У%"Ǜ��P;�) T�}�����Ȋ�u� �l r~K�i�A+W��C&�/f�|,y�����x���M����|���^)w�z]%�|����aKR��Um�'
�P�D�A�<���$����>jI����~�O �x%��e��%_����#C�,�'�q�a�G�����
<'�E8����9t��8Y��iUޙ%%��ߖ����ο�'��Y��ñ�za}2;��(��3�Ġ�y +��?:���,7B;��@M��MЉ�ȊݺMu�t{kDJ����p��8nP�6�V�<����f����G�|hғt�����5�oH?�y}��Ɨ����#�}��zc��j]�����@�}�}�[,ʜT��a���m�Ŏqu%�`�gJ�!��{�T������ql(�^.(r�V��&M�9���h��t�Y�'Ƈ�C+ڢ)Q�2t��+x\��*�&M0��� ��V'K9�ț����#�1A�o��*�FC14WSVڑ�{��J����l1m������精�=J�s!���*���&\.񗤎gq�5Z���*"��(݌Oy�5g6C�v?IW��%�7Oj~A�+� g|�1k�HΓ�����E���g����l5���|�'b���ǚ�V�疔�����;�*��vP�0=Q��$�NOe�� ��j(�JM��� �J"�Q�z�!A.��gy�s��r��bGtS�+��͢4�
�ުȝ�S�T���:�|�������_���?PDd�_��A�&f�Bp��L�A|�(Z���@j��[��
�C1�Ǌ)L�b5�l^?bo����֝֡X�ǅ�J�:�� �B�*�\gx�Uu =K�睐	m��R�D�ms{�y��%�wgd0�Jq�w�n?�޳�q��=��\GL�F�P%-L ��9�����9�Z��������):ڊ
�*w�Qŏ��G[o��z��F�#gܿrT�.=�������g{%��E�,�j�p셇���@2ow��4��Zÿ��3��X�塭�1�h�0ܜBӄ��n������6�[�c`�qÜ�H��R&^�Mt��IA�֬��Ŵ��؁�*��#��Λȥ|4̌ϤzMr�0����`"L�r�v����wG䳗���Gd5ĺo���v|g�����Z���ۯ���C+X?�*�����ǑSW��vd����Q[�=!/J��Kġ��b��S/��:-^��Q�5V���RH�/s��}�jeőbB5�݆�+��ծ��/w	��M�D�?r[*�����
�vg/h�{���SI\�ک#<��ε�l�������wF��_���!O��3q'ddixP[F�;�����[m��׆�L������Z��ùA��q�]�2d�1[�t���yB<���0�T�fʂ֊uU�����:���o=�۪Z�Kch�@w����H��Ÿ��F~rɑo��6�1p�,�m
ӭ�a;�[L.�k��!�$>@�b���S�+�G�ٹL,��M]_8D��C�v��� �np���3� L2��G�}��}�ޤȻL�i�·���:���MTd(ʴ��6��]�^��n�����d]�)��6��4%���¥A�Z�tb���I���T� Js�;���kɨ|P=p,�0��U���u_���X��]�$�tg�S��.�\��A��YF��(�y�[T��hQl\���2_	O׈��*#^P�S�D p� 2��К�M:�ʣ�[i �i
��t+5q�O=���	��<�����u�l�g���Zq�:�� ����� m�`�v9L4�rf��8nYģ�B�qd���L:q��mu�F�S�I���Qam9�� `�J>u������ _b���2{�DL� Z���HH"�lx�/-��ܪ��H)�i� ;3l��[����<^DƉmҟ�
7o�����m{�=u�v�!�p��v*��K��D������L�sk��cI@���ȯ�$U9.��كμ5�$-p6�P�'�@N��D��:)�Jc~=/�wqަ@�T!7V�P_���M��Q�4��\�U��Ҙ��L�>���$DW<�t|k3]���S��d�)M�.�����溶�9�/�e��
\ɬA��X��zsD�ʤ[�S��/�2�WKK��ϖ_
��'��H�&D�o��1�\�[��42��c}�b�%�3��/F������Ok���:)G���f0��S��Xeg f��|���cPD
y��_��WJ�5����_�{e������%���)�'� �U��m��9���2$ ��SJ�0�ğ���b$2�D�P�ٚ|3�
����(Zw�̿l
� p���AM��8�H5=�d���)z�/q���6
��_XV�5���֟6�{�I��+?���;1��R;8>�D8�j0� �bX�$ۏ���"��N�ŷ��`�qD͠��cё�U/�K�⒊��̛�%�F=gi2�N>��4|����K�|�Ds�3�<��l��2xo�[��]y�N���o�*k�Q K3�AX�H��6b7�ۆUv�![������F��oL@.e�]�s�����2Z�H��bMa0�(�cO��fF�In#�S�j��ŏ�U��3X"����o}0�V�N^j�������>��F����h��ʉ�Lb�VN��7p�ܼס��Ўp���N4\�#�:ֱ4� �fkIv&�[��)�3g�P	�+�p1p`����OHd�8�^�����z.ĦEQ��RF�~��V<͹<~R�V�f�emȀ�o9���)��jG
�/r�!�u�R�@���^y�T�)[���n>���D�<�2)������3�H�2���F���	v���5����#ג[�7�w���]�P��B�{YYUC7�XM�\�|���.a`��Tk�_�w����1@ۜ/�);����M΅1㵟�\������$���
>�1r�s%��$�C����2��R���l�@H\r^�E�C�kAVo��VP{2ӑ�70�t��NQW������b�*9urtG���o�� g��4o����:xwP`f��gg��Jw%B���6�|?�Z�#W'b��>��<��[�� d��/%��Y_�$vr�xK
�
H��`�QB��m�wq��G@��� ��{Ⱦ��HA�n�G+,!�Bs�"�)�»�f���T5Wj��3�6+�Ë�!�.���t�9��:�F��!�`f6��fa숷q��7�ş�~�bw���-�ud^�?����a�wl4�*�k�sZ��Z�	%��g�z�%���6���_�z_�l%��IS����rZ���`����{�vn���>U:8�]Z��պ��x�5t��^!Y&^;A�A٭lǾ��a�։U9����ը��ԟ�����]U��0OEb���xɌ"�/ ��������W����p���.�ΏH4C��o����0%��?�Ӟ�Đ����z 6C�?�C2>��H�R�_�陻�TZm��4�e���SG1sa����1Ɯ���j�5Ќ����βG�TU༛F�j	�t a$]""�_oX���j��y�.U�oiM�
�,ͣS�X�kb�T8�;�]'�e��@���O�hP��6��?.�@�z�8�3���� r��k�����`W}6�V�fu|�	{�7�Vf��vBƠ�<&]�i/��]�u�KW�Θ#��Z�n`"�yr�!�.m��ɖFE�hHDGr7a�ѕ>��%�ǢF��7h�_��	3��@zQ"�b�ƌgi!j0Ź���WE���Bᘊ�=$�l~Ҝ�T��x���e�ӥp����YXO��fB��QzL�m���u�/9�F���&��$��~�}J x��wgk�po=���N�_��X�
�Ȥ��>B05��S�����fn:� r�2����B3���\2)�mB�LsaCeG@Җ��3�tG�ղ�'Lb�M�{���������O8���u;w�F�4إ��1��^�z�|��.�jm��/\����ׇa�����>,�L��s[��L礓[w�m��Xx)C,�|��B{��3Ꙛ�L>k۰��L"�֤�!�g5b���C���P����C�N�^i�e����k{��5����CR�UW��[�<Pe;��p�vc����x�q+,�A�`��dB��>���>G��.�Vj��3]�r�(L�`t�)����6ۊ�8YS��]D\�:2z��XEYU�	nb\���9m��9 ��º��Ś�y���jr5��Y���ꦬ���{{4�����2-�D�$a�__ٷ��v��0`��.]���+�$����w�� L���?�KV��i���H��`X�P�I+0Z����F~l�|���HD�����L�n{�Xv�g%v�6"uj�3/�$���������.�@��G%�2�J���jpz�h�2V?���G���+��fV��#�E�xx.~�9��>��,�Yڏ��H�����D��w���C��"�}�<�k$h�k&��5��/$(=��S��{�z6eْ�E�+��@��rOg1�b�#�&�dG�v*�s�\5ˑ����hb�r`B���l'~OIg��Yf��]:8�y6S����8�R�s�./�Ro�$�+�!��)1>��:��&���GW��ݿ���]~6�;�&�27Hˉ[Cp3�,��x����[�]�?������C`��6rTX��G��O��d�V�>��>����3��aʶ��"<!�QB\�!0�:E!s�VD+���j�v��,N1��i��ۺ��Z<J��*�B��ÿ�]3�Į�7n�V�"˂��>�����Ō삅�=^����.^�M�IF��	`,���<B���� �O�E�ޝ#6c��pg��܉%��`��nc��>�Ɨ��$Ȓ�N�h���*lAC�%+���+��s�Ko�-D�p9�F� #6_8#��~���k[���n��z;��4���p�&	�a`�"Yw	�A}E��rǚ(���̆PK����u�*�4�.2��i�p�jt�4"�&k(ߧn"�,H�������Z0�Ң�~a�`�*�-��*���%�d8����{i��~�J�����dw\{�X��B�Ǚ�t��b��`j�P(�@�m��m�]�ȵI0/���VZ�[��zZ�r �-�����T���`+8�Ğ�P(�ٟ�R�����w�L��JPߴ��
�
��5@i�����E|퐾�5����F�5�Y�"ܼ�х���?�-
�u�t@S�%�±yoUx�u
���e�>4����˾x�����&�8��eB�C3��?���L̶�h1�=����ڎ#LY��dYЅtz���~�8�4�r�Ad��ƾ����/�D=���m�͓Ok�+
�M3����4����+?�'z�A�7����+�p�gT�]��/B� �73Ծb>s�&�z͘_�S�vg٤��9��C�PU���IHh�t}��4�$Q����Tf$�h�~z��[��l	)�OBc.q��/^9���|�p~���"�hw�!a&�Q[x�s�yM��]}�M .�i��O͚9N��ލ�j)}����z�s�"���M��	`�����p[%������ix��iȾ�ǽz� �aAh�w��l@�Fl���
\Τ�S֭~����Rl!�F�}��<�h%5���P"�O�I��!KN�g��qL
,-�^��g�TD>�g���,��>j6]x��<�.�h��lN7���*<^!悔܊7�� �	�,pA�cۆ��e(��l���VvL� �Ѳ�"J@ �p�mGa-#�������ё��t�I�\�ٷ��e9��G�Fħ��\�o�%Q֖B�[��O�i�nK�OE�ja�u+xcJ��c�/��l��j9H���z�*(�>_�a��hȺ�s�X7h #-;Ѧ:X���E@ԫ�H0g����B�Py-�io1?	,⋂j\H�y]E/�����D���$���+�fƮ��9�u�r�p*�S�jtj�lb�њT��')�5v�J��ǰ;� �����J�W��棤�;�|>F�y(����KT�M���la����U¸�{�G��� ��ƞL�d����ܠ@?��x"W:jk;_e3��b���'����ƻ&�@���wP�g'=���G�P���!�՚�lJh_��L��!hJ1�_L*׌]�/쨥�B�f��`]w9%���$��?�%-p5�T(�ю.Jۚl��a��@=z�_�#�IKL��B�'r�72���+�?�}�R���/oۇ��B�C��p���w8eT­���wN˓���^H�B����~Cz�03f�5�{��C�G���^H�[���YՀ��g���#�a�D�|D*������\գAB��ei����:�xI ������s�n��ZI�.&�`�^�����}���&�xk_A˲�WfɊA}^��-�p#��B;�{X������/�>x���/F�"]N�����O:!V�}�@�/�{gT����s]��?Hss�J���ru��}�d�z���:ٔM�%�m�bHSx��m�� ��U(�ߞ��e��p���财��~D�=�9�ة{h�V��L�3�0���J_�����U�6���)!�]�����l���1_�gǄ��|/�,67��Cu���D-ݪc��o��HQ#k�KP�d��g�|��Д07�9KU��T�8���2�� ���7:�k���"�4~H\r�k��������A-((�="5R�(Z��EH��-t��6�G|O�3��?��u4�LC/�k������T͕Q����E!�?M���I�.�}s���k*����Q�g3�y0u$�2�^V?@3�1JI��kuї��a��4I`�L�S1�����]�뙯�3� *��7�L���D��%
�}�o��E����%�L��5�o��COj��/�f>�n�Q
f-�5ޘ�juc���S� ��g�"�dz��`���A��[�NW� �_0�x�-�5�? &����	����T�w����d޼�,�ח:��a���<���_+�6�.�_H+�R��VR<�?�����a��8�T�o`ɕE��$��X�
=3��ϻ�_'�J^�Ю��(��Fts���=)��ƎK,o�*�fAMՃ�֚�q��6��������Ԩ~�*X?�c=[]x&�N�>³W�"�qbW�@�sti���ٯ�o�ad�E�����o� �12��L�+�g��'�`�%���1�K�5��ƙC;{�V�cң��U�H<�zf�(<�,���ю*#o~�Hp�ʘ[�V��8�F�農,K�d����riN������)]���B/�&)Z���"P�8�}�"�ȓ�(�7�Ĥ�iY?�W�5�ٟ�1�^81_+s4����dL�a�����Vp�����Ao)��﹣�Rr��!����ҩ� ���9ϗv��@;��Q��S��@�_��8@p1{%'�J-S�n�7P���Ŋۖb�m�d����p(��y5g�S�����v�7��om����7MS�a13y*���B�F�AK��{BO@��pE��[>�"�i�0����GU�h�_#U�Mt+:�!G;�3�w�r��-~�7��S����F��Y��)AOV3J9��Z�JG�ht���wP�������s���2V��q4>su�Z*|�tMV�o��o	�?d�/���4�����w�ZQWP�=���#4޵�t�鲚�(�]���=�mO��9)q��R��S�BӋP�Mѯ���������ʁŜS�	�E�#�K�L�0�*��V�)�lNTO�׈��)U݋��H$h�9��je8EW��6��9Ϛk��$���,L�=f�9��WK�T:]K7 h[V����R[����m��;~������|Pɿ��";܏�<	���1h��=\Wa3j��вd��s�N�9��CR>;9x��X�f6�� ��B�a�V�R'?�Kz��F6m�Z�؟Cp:��k���ڒ�!i{9�Tc'n��F�!݄8%.6��,�|���.��9�CLJ�'ʽw���
��8OS�Q���5�l�%_9iw.�h%v�Kx��|�Ǔ��ȏ�j���_��@�~9������U�:˒{哚�3��,\)f��@^�P��.]�N���M0.�����B$�3&�U���V{�1	��'y"ձE���$KT��Q�	���2Y�7K���J��&���R�Z��a�(lг����VOp'L�d�Q.R#i�߹���3i�лɩ�7���f�j��ՠ�$5�C�%ʯ�����z��&��� �X�
;h�C�@���N���#�����/��q����(�C��:�`	i���p�8]*A�֧\���\E����4Pz@˖,�}9��L^
Qp,�G���S�F����%��B��}V�JK���X����Y���iq�Y��E�nY34>�0U�y� ��DP)KQ󣭴G�oNI�U�%]w�N�N�p-_��^-?����� 7K1�8ұ\���9���vN��<m1���1V��gR�!?�nJ�/�΄ί�\���Q4G�yeET:;��~tzZ�,j8�g?]20yԴT�LL�;�d!�~�5�$g�~��K�^�@>�,��q�1R�SAi�TL����`ᪿ��T�S��շ7�zD;+�{����Q�J{���z���Ku�c�����c5ub���C����<ס�ɢ�Y���En
��h���1�r��^	������%�0ƻ�39�9A��s���RTn���9�YJSI���9���>ۢJ���2���r[��
1O�`�75�пl+o�ң�w܄���
�+^(�����i�p9�9z�Jb8a&��b�#�`��:�w��=�v<m,����&��X�V���M3
I|�}�@?��*=��=���c�vB窚� ���\��Ǌ�$	^V���AA�S�l�����ԙ��%�T�!�0���{q��p_Bc�ŀ��װe�'�����n��	ty����醢�u���@��C���H�.�;�!�'%���}� ��`jl��."�b\�~9���;��{=LM)Dt���
v!J�ƛʱ�t(��ԟ}�G��<����E��Ax�-�R$z���s盯Zs��}nɽ'����ZSR!W�~��5�1B�^�'�7t���B��9�'ܓ0~�P�S7�q&muZ,����c^��N�]�2���|�>	U�*�8���.maؤٛׯ}��H`w(�����3�N���*�F������w`)M5�xA��	e, ë�p�tj�VYH�Fm]�X|J%�����C]�PU�t�T ��������0Mϓ��]Y��|�B9��z<���W��b�x�R)�����i#	�G���Æ<�1Ș�:����:�����v��`�L���r���l�GM�B���b_�x�e��̮:B?���(�Hl�� �ҵ�� q����=76f�.�WP�ƥ��{�P��M[�4k�ǝ�:x�.Mԓmx<ϼ��D覓�fwn�7�<,�,������;oyO�P�9b��-���4��2��0�\�G�z��c���I�oi��!?m��p��|/�f��Fyv���@�Ҳ�e���؟�wAL���G
l7������}e�5�
�� )�eD�8����C��4]d;���OY<@`��A�qn;���6�"�n`WE,=��	��_ؐ'�����o}������t�����)�����dbfB%���5�-A��S�+8D���z��	�g� x��R����)��԰��v�d"Ib��W��8gg&�=2j2�.��B�=7�6�D�O��e."J�"��v�(�U=#�7���f�ֿ�h������D�ci�j��Dy��Q�'�+C��f�:�����(���*��-'��dby/-�.�3��q�T�~�Q�u9ˢG.���o<�fcZym�����36�?t�����.��3����)��L��?�뛱q���.�e��=�PJB�2�K��4�|&�	(��Sr%�7�O+�)^�����L����ݟ��9~�Rnr�d��ywo������K}���q��j���V^q��}��S���9�ݖ�)Z�p��Z4ej�D�!�h = �a��&�.����2lۛ�0�_e`�w�R�F�}�7��c�oc-9Ͼ9�}��a��Sf%���8����-6�����%L����z/��NJ�/���~4�]��ܐ���ڏ��G�q�Y  ivz��\�v"�zW5a���A�!]M��b�ysI��P$��g��V���	]����,��-��6�p]^�����G�߇=]��lJzN�Ol�r��4�.�E�'.B
̝��|��Ĭ�_�C[�M�hg�N�C)�[Ԫ����Ƣ�b�2E8��Y�����(h�.�H�W�C���]��^)���_���u�����J�H`N�|X_g
��DE	��*WO���M��S��/`Ҫ]+(�<)�r}�+��+2r�q,Q���k�Ԅ;���;�x2����9�q/>ej����<�9d_~�<-%Rܗ{�o���s~���i�s�6�s7�&R�8&���s2�S�p�)Υ��6�f�{�o?����R�Fv��SJ���l؋]q�VP�	}�@KM�y���
�J͢é��1�t�ޯO�� �s�',������M]����������9���?mq[w��V(��@� ��b5�z�<� i���O�-6;��#�A���5b��6P|ק ����/��6Y�+��i�@yL|(7��м>E&K�8���M	6O��;\�i���9f�S���e�D`��3(��y4#�H(I��!�Z΂Ȍ}Urd�Hs����~c��q:�W�G�]���lR�Rv�.�y�ϝ�.�;}֫��� <V���B0s�?�G�r����b9��.��UpD�mI��ꤾ�1�؁)��a�q[)F���yۚ�� �3n!�P�p�X�k��0n���������3<Kv��2Q&/;�O�ӊq�#�E���`��T��f�N㎞�5�0��n�EU���2ES�n3r�R_�hюXR���7���y07�\h?ƚ/��
gp��$�%&�[�Ԓfja����b
��5/Y���o�Mw>��A���(���3;�#}�U�2�'^��u��E�U4Ϳ���{@��#>݆�<;&u�_���p`W;� +5W�)����}�<�om=b�,��l��8�OL'�ɼ�6�X�i,`Z��r� �sjS�X(�0���ZD���7�E;�U�v[�vO������"�֋�@�`��T�Hޏ�h0��؛��A�݁QnV��:�jd|M6	�nO���9�OP�+������2y�$C.d���A�&OS_��6���a�O5��+*Q$vrZ5ba��D�'�4A��]�e��ظ�ۗ�b�6�q9��Q�\����$��4d��>�a-�o��@�G�6��@�5�k$���|QP�,�r����T����u�h]�a�mŊCYUv\u�.i�����{���Q2>}���8�a�[t5q+�N7{$c9�:���F<�df�5�Pfjo�,j|�kV�1�
ŵ[	�&ށܶ�V(�D���F�
JQ��\+�v���u,����2�IN;.��@�(�=�~��Y,&ǻ@��󘽬�A��D�
��>�h<����=�:9(2��b����Bnh�?�[�~)��y�Öb��X�"U�CN�V�ob�ݺ4�o����&lؑ�t����'��0P��:A��+��8A�S�!x	bɦ���1K6�����z"i!ko����׷&D\[�1ۑ��Mc���2������FI��_��@�ն�(�jg���[�]��X��er�ݗR�jJ/M��e>z�K~"�/�rm+cE��tW�O�+�lC�w�	��1Y[�d��LG D6�lg��\�Я���0� $7/��;���;�$w�Q��oޚ�E�+�X͵���Dw]0�-�ѷ���R����Lk����ÞP{*=�s��JV��o���B�Ir�&cVf�F@���/Qa�����*M�q0,D��?��BDnv��>sh̼\��k�5"�_�C��~�],� �y�j��Gd���}�y���:	Ibx2��2 d	��nu���BgH:ώ{����_�vX��,u﷍�Ե���n$��Oz����o>�W(���/�Q}�3�爊�B~���5b����x�cԸZ)9�I,��݄m�~�F��m�����=h����>Rz�.~�=ZV�L��WN�P\i���c,`��4b��[��V��I�����c>�g��E�/���3�Vj�
�Z3�.yeHS�L��t	�RY���:G��.�v��M�$J3ɯ�P��]2ˀ- ��!�+����� �~M����(D���L��d�x�A��J�9�����r��w�b��m��yx{D�['4V���������Ӓ�]T��-�sǔ~
��!&K�4�Z)V3��mTd_ƳdL8���m�|	���22���In�S����Y�?���Iᳱ$� ��(FJ�KZ�a��Gzˑ�h7엌����V���~M�,*��������n5���ǺL�5]a�����@VF�*a�Gt8x{Yv��?���
�9�Ej^7ȑXp�W"_��SuT{B+�$ 2��^����&J����&���8ͤ%��e��i��8����CJ$h4��-F�Ӻ����J��V��;2n���0wb%�t�A�܏K�BV�p+��y���O��{���u�V�x�9����D����ͷ*XX�o�j���'��5����rǂ)��eGՊ	4o��RQ�i��T����z9�G������I8��ވ����F��n�p���i��z���kO��q!����o��B]�Q�1��ʀ���Y�E���Ô��	�j$'U����B�%���{_��?!&�L����8��ϼ�8��v>�}�a�e�0��ew��m�
/4�(w�I�ԋ� �����<����n��7�î_إ	=z��I�0�G����9����'�6�?�����Bf-��,���b���O�g�t�۵��<w��-���M�ö��J����"Zx�-_�[���P���w�kv(M��ʥR0��5�3�W���]�+`i~�2�Q��2Dr��^-��"!v^b*`A�#)���>J�7"���r��d"���__&|x5{����� ���N���1�V1s��X�RN���4��s{Z�N>'�jX�#��L&=Š���=l�ϋ��jl�d��ֹ�L1 ~�*�m?��N�����΃����&��)���TO�j�w5O��4�w�_�|����� sD�fI����_K��HJ����&��mi�N +��G�x����ʟ�m��?ퟪR��vG��+�\u����2���l9"O�l����ך��O&��� 9?/�d���>����X-V�׬a�(�~W�F7�k��n���|ع��/
C���$~��N���ۖ�/���<�y��pԁ�� (Y�-��W�����sM�'���WYa�=�y�qd��u, Jޕ�}��C�d��]�l�$A_J���;�y5 ���`��H���pz#�S�W��WbU5*����H{�K:��۪MkuVR�:F&_�! N��'9Ӄ!^8U�����F_H.�v&i5�(�|���-o%8kt;R��=	>V��ho�$uhHWAd*3yd�DK��?�|T!#��Y'�#�΢N���?����
ù�.n����*1��q�J�P8�#4�k�+?�!b�X`O0+�G����E�j���i!�K-V����ɶ��)��

��m��І%���*M�	!�-P82�����X����5${��*?�r}c��W�	l�0��!Á<@�P�t��L$:qɉ�{�`j2t�� x%<��쪪93mZ��Hj����LØ8D�Z�#�-����)+B�So��(2����!\{��-���k٧��ԤY��!H���$of���&�����Z��ᱚ8nuX�`D����,����1n�hD}�p<6Ŧk���Gܪ� |������6;�?����ˏ)��(��A�o/R���鬱��4_�:L��b�gzX-���dC�w�"��l�̥�y'�_?�i#B�!��-ڤ�	�=�̊�&���������OP#:d�(�[�PAV�����V��M
°r�<�R7Y<欂� ��\'�U�k�V$���
�.B�69�C}��U
�4.�7����2�Q�4+5���Pit�6���FUG{�1�T�xYA�aЫ=v`L7b�a/_O���@e���* �>Da��ޮ�0�|p��K(5��_3������1���c��Ŗ.ρ��|W�"ǣ6�LmaͦQ��I"�m=EA��[*卜���Y�:�_Zޓ3�'���B2_%�+����'Hܲ�C�S�����>0�:�$N0I��c��D���9}�7����>�)u �u������lѫ6��0~�җ���_Vg�#�{�K�G����\]����<�����)����;q�F�娒Ҵ����J��E�GH�m�,��,�����@�L�>��C2;��P��� ��X�b|Gz�0��Y&򴤏G��,K�ߢ�3�N� ^T�L��"�u�����+͏x2�BTs 9_�D2��Ph^��+�zB~�3Cj�!��4DЬ*r@1�{p8�t���xgg���J�p��mr,��8�!B��(�\��K��*r+�zB�
«)�Zh��M�.��;�\R�|j_�6B� P�����;�]zB���|  {1�O�\���M�92TI�<=������芻���/N�C�5ߢ�� �~
tuPђA5��� N�f&�,�D��7�(��x�&�'�b(�����=P~�q*��5{[�\���"r춓�D���G��Ӧ��e�@&��0�H�%2j����Eú��O�`�fm�-�<|8*�cZ��k^8����\�i�wۭu���w�wGr6^�}��6�n�i�/�*^o��sf4ŭh��J��>^��J#�>^�&#�+;.�;�[ҺL�H䰔;xvٰ�(�i�f�ܹ��Fs�c'o���x��hb~~�Ƚ���ȧp���pR��]���eD��l��:p��`��Ѓ�}������2��!���/�ÃX��g/��������L><{}�}?=�?�?򂪱����G���ٍb�+)^��g�mo��k>u��]��W�0~Dw �ImB�f��N��d��GP�Ei�}ۓ�)R��
U(��-��2\hH����]e"�#3@���-��,__�!ݪ�%+2�S}/�o���)���a��\g�V�|� d��W�i�F��&m (t���R;�@��OE/����
���$ø�bP�հ~zq��aF!��63�߬��K}���\l�CG=t�ŗ�!�%B���V>����'����P���/��v�ߤ��4�Z�C��q�H���bY9Q{��j�ހ�$p��������"�T��R/�.^a��˕�L�ɚ⌭��ț��3zk�	~��Q��9���3JXA��(4g��9��}T�v��	�}�N�Ũ_1V����C&TL�Up�x�.��4Z8�xE|���:��MA�W&�>w���>����e��Q�XǕ�����
at�p��q�v���늹�D���"�b����Q;	V�!�p���f����p�<�*���s�-��%1z���;���"�q���O��
>Ez&Y��uɱ��lrƺ��.�+[���(Q�|�V�s��G:��w��R�rD�Ě����d�k�7y�-4��h��JW^��P�""gqt�9j�h�n�i�9ʄ��3����u���/�d���RW�ޑ��I���a6NL;D��Ƭ�vg0
t��˧"�d^r��DVj���F����{ʘ)�����Q��lA�����{5��n9��V��c���T}�?Ĩ8
�G�p׵c�e�y
�@W�dW$z<�,o*T
�����Ȗk���ˉw�>�f��^D���W�h�y�L;�hga�`8:�)�e��m%-�R����H�9ڂ��F��������i}'���Y��J�Hj��(þu��)�o��Ǟ�M/�|˥|j�n������0_Y�Q��coC�;u�;�
�HE�H �-w��bWg@�1|k��+�X��,���N��5o�[��A���ۙ�ǰ��6�6�Y5��|���=��1��_���x��B���$�;KA;}�f�>� '7��c�<��5�s GĹ>��1�����+�
��웕�>bZr!w����{�fW�H �@��W
8HK�������\��^�ҥ��W�%�b�/���֒e��/2�g�1�y/��>�O�:W�֍)y�f���qp�J��ͨ=�S��"�/���Z�Q�t�g��NRjB/H.aUz'�D'�1U�寜b��+T�÷�H��u��J�9����6V�h����%'���v��4MY�xJ�'~V��q`�� r�&%��+���6+-��c�섎k��lr��&ʹ9v��|��o�w2rc"a?�Q�?����|�ܶ��앟�Go�ݘS?��gpt�C��NP8rv�E3���:'!�6�,�C"�\@��W�މ�j"�Rt.nL��Ὥ�x=�?.p.�Fb����9|�L���&4�r�j�j~���њ«5T��0�`&��e�;�˴^,�����[14Ǔv7�S��Ň$A%KV_�����~Ź�,X|�4q((ow�'��Lm0rrx����~��V�6+��M �)��U�W����lu�[����QR�Px]!�^������������Au��Ԅ�#kf��L�.>>+�X�v�m���:B|���#%�P�ѯ�G����g���Ty���?@��խq�a��h����}�|����FzU�m䕽�9��an�	�{���q�u���@�<",Hȅ��b8�G����\��`.�(b�x�Ŝ8j;����X������
F@s�G+n�����ռ�cd�����[���d($_SS�^-n�gghr��Q�/0;Qr�*)E����>�<G���.٪	�OZO*�dt@�E�_�g8�������0����܈�
E]�Դm]~�ٮ��u��d\��#S��9���Z �iŠ!>j�\������
쾰��΢�p�щ��I������NĨ>'�`�^���0��4�9؛C6��M�����O��b�a�'�"H$E���Փ
�W�'��T�K��.��?7�Ʀ�{�1rK��v�x�mPib�hT�,�֦v�A�>����=��J����v���Q�Ux�E�mP"e%�9��A1�η�u�/���3�N���gJ��������;Şg�P1y9u�b�-P� a^�F^�&����D�Œv��ﭼ\����ȅw�!���z�S��|bi�3~is�*�n�n���v�&^��5�m�P��Vݚ*/r$�}9�r�Dr�fe^����c�^�=���
X/j*Q=삤-��H��b��2����smu4�/�˙K�t�,��y�`��_*�8������܄I���T�3���-��{�5��0�qk���X��' +NY�Hi�|� /(�)9�]��f����F�1_ŝ[�o�>37�x;w���fh�O��s&+�`3�\o�޼�-�Q�C��_����G�i�`&A5��E��<�K�D�ap���9	��~�[,�L4��/�YC�98�v#�_��/i������2�-<-�2����i�i�ܹ67$�MZ�#ށ���nu8�Qw���cp��\�dWq��{�C�@���/���1� t�^�d��T�b�E�f��z�.ѝ��.s��Ǔ��e�&�%>�$�=E��B�	���qq��%H�$)8m��h�p26گ�vL�X/��V"�n4�n�}�V�< �IkW~��c�n�_���zQf���'�w��,ܗv�t/F�"�cn�^#���(��2$�V���rf�����^gl<���a�J�k"-�3�)_	��F/~�c�6�'�w���J��پ� ~4��:�끌]���]Ѓ��9�|q�y��^��c��U���rߜ	�A�mg2�k5��pkl��Wa=�8?g[���b.��|��%�؊>wT�?w�U̦�����L����Mg�Ys�٤�VF;pw�Y��.��yù�U�q�CJ�*�5l&`2���m\�˹���=_\&�h!E�X�,W���#��C��fܞ����H�WIt��rQG ����5�������AUd?���r��������*/���<_�z�]Q�5%�_gj�]�C ���ŇМF`UD�I}+�x+lWZ��=UX�~��0�@�S���#�r���Q[�0�w�6�_$��%��PDڝm$�`�uҜf*����FL��|\櫚N?ˇ��	)�+�	�;)®���3R-�v�֘��
�u�2������}π ��Tev��G}���*�Gd99]�l�@χ�N���_.P�L��B0~�-z .1[��#Oq'�IY�}+���o���=A>#�i�{�����On��ie軞��J�`h��d�~�����ʌ;�����͙���}��0.$���U�Q��������L�8 �x��$O�;����ݔ�0A�BN�O!�r6�$�Lj6{�­��3�i�>�Vg��j��m�G��C�#��mEA6�ǜ�j�OV�p�mL9"Y��O��� q�O �(P����X8eq�3�p�N�	�
�V�lj���7D�zr�� /����� =�'b��1�~�X�g�A'n�\Du��Ԉ�Eŋ����*a�)�B�z��٤�7C���]O%d�2����<�U�C�;�J֯$��M�ɖ����J�G�ƱG�=\�n�F�_��1wA��CM,� ���2�,����)�`I?�ne-	Z�a�i	7������������MD�{�B;׵>#I���I�z`��'��l�e�B����ޯ��:�HF��m���ա+�Y��֯�M�1�V6u��S#�4 �}[r�X��;���#�闋̽�T��U3�3�*ȁ�z�~�Aj���v�̜z�
��I�F*�������[�iIy���.y���&� Tb����ٽF�]��z����R�Й��0�!"j�0�R�ͩ� $c)xI�Rm7�T*M�1�5����xu�4��q=S�^��j����.n�&.>de1�}�������4K]M�ګ�8l�L�Quu�^���!����2�wI�0qNrud�I62���8 ���(Ȗ��K�'eAX���lG��c��c>���&�f�����|�2�`	ބ��W����T���x�C2:h'�ʅ �~&�vE�1��#F ��a��"�8'�xYz�Y�{!��\	��u������p��xz�IC�1wb�V}L���v5� mW�.`G.��M�m��?Ë���m_��Q#�%:��Zv}`��mG������l�F'����a�����ʙ���[-|�����~D�=�q,������T�
