��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0x��lQ�އo� ,�,.��GtZ�.	���@�'��(��uL�X��$z*�b�H���vݹ���]���z��b�{�O�w�.�[�i�go�(%� �]�Z��hp«鐣 ����~�bp���E�+м%��0ŭ
���8NM���$����+�f@�I�l��M�A_�᭼�]ƾ�$�|Y����|��A�C0C3%��OT�'~��!��|R��QF�B�U�' 7�b�?w�!��|�'5�)�lL�����{S2�)�>� ��QV�,�D�2�/��h�69�6ܟ�d�Ϋ	-20��%�F�, :���)͔df}4��+�p�O�V�$���E�|&!��l��sN<��lS����n�J2Ƿ�sK��۽v�s����D/Ӹ}�\&Ϛ�S�M��%Ta��0rG�������DNʓ-ݯ��y�S%̓���%B.-8GQ{M��rΊ?٠v��<����!8�Ȃ��7��v"�zq1=����p)r��`q:ڑ��b1K�l�1]<��.��J�C�����ɴ��b/wSP��N���p��EHvD���<Jlk0k[�p�5N+���`����W.�-��$���1��Gh�D����MR��Ì�$	{HC�^ ���F�2JA¬���0�QE,�Ҹb���*��g�s��gQ 	�/�R�	�N����W��s�cZ��<�)�}�DN�> �Ϯ ���]@��<r��`_��2�D�JP��4���)UUԐ�� +F����Ne�p�#�� N����0 �@�ά�倧Fr�c�F�%�l���K��6e<�?�C�aT���X��4�+t,I�e�:3@�K�2P���,��Y��Ⱦ��˕p�ע){ ��|���}�¢�1s���G'�֞��^\�W9��Y���"��a324ka*�)���R.����3�,ɩ9ﾌ@p�o�%�B�zy$E ,��;Я��¼^�d-�����B�j�:�$�Xc0$�W��[P���(ǡ�O�q[���6O�s9�o�Mo�[��H�y�d��$�
O�vţ�ʩl�����8M���};���V�k�����|@�-���Y���6�_s@A���ʉk�&�U�����*m��4��������}�d'+Wb����R*>(�����hs��,u�����ƛ�����/��V��qH�q]`;�^�^@��;�aB��ݯb�����L�v-a���B(��0u�3C��0UEH�V�S;���S�Xd�|D�bI��7��d�J�E�/�<`1^O��(��f5Cy<n/-A��V@��d�}��j�dds:�{�$������Ǿ���S[߻������Os�7"��|�`�J�Ʉޭ��s�*��xm�Yz��@����{ @�`\���=�0߃�ֲ)��4<(Cs.�(
,��ft��0�X!�&���6%X��������Mщ�L��v0��'�������k�jpy�����EBX��ey{_��Kڄ)��ԯ�=�,fl�X-� �ࣷ�e�R����`DpO����Xڻ�&k��̎7�|�|OF�7{>S7W-�PPzѢ ��4ŧD�%a�]�������g7��Z9�NP(]�x҈d���[�?�N���{�ō����+��@�x��R2��ƽ��#�: Q�+�������$��l�e|ے+��M+��(/�N�O����"���8)�n�q_�#;�(�0T���`*�J�
�P,�
����-�b��j���N�"�8 8��q�)r�n�8|��F�J��((�7�ɺDU�T6n LM�Ĭ�8�'�fos��v�:,QۣuZ(
�L���Ҝ�C�F�ʻ�+���?C���V�4��7��H�~��uKq����d���TՁ,=tp��݂6x"��u���,�����`T�8|��p��
d]��w̨�1`��w���O�����8�p����ktޥR:���\L|��wsI�<ΫY�T�q�l)�0��t����k$�{�<�,�8m���n�yk�����p�T@�XU��&��_Ь��	k�2LMl��弘���Ik<zӣ�A>��9.ϛK�J�z�8H��h/��-�@���aq��ZJ���B��(�Ҳ�G�΀��g؞s��nԈv,j!��r&s�Gw�O����iP�y'��sM)x���ui��[�Gp���^�CWq�Q���tߗ��yԓ�o-qB� ��E�To��ʧTIz�Λ�[n"9�X��$0z�6$&�Z�]?��cok����బ,���<d[��Ta7���z�����3�R��Y���*��,8Br��J۲��&�6���tp�?B�"C达�&l��p{o��U���5��QS1^���I����AULF� ��ZD��3q��?qt�0xSgtoF�p��WJAC:��x�3�$���.5�t
lz��=#Y}��4�Ǿ<.�!�;��C���v�Z>;��1�O#��	��30j�O7ZF��%� �)4�S9�P�F6Gђ�I3\	������W�4�=��fZ�n	4�4���2�L\�I݊�Gy�]˥Ȅq�o���5������i?��l��`i}�8���s���ddx@�|P�ʒp
]��l�?0���}��yiD�\/
�u&��{��R�;,)Yz��Jf�D=%�>p�+D�d&N�#�s%�"�09��[����/�9^�-}�~��k>�JM��oA]ghA� �:�����+�=��+<ò��u�~K���݌���Áp���	�3��; ����$PyY.�=��{&h��X*��0j�]T�	���YGD�ѷ��Y󾫹�ܞ!
���U��L;m�Y�AJ�(J���M���㴕����W�!M�fS�d��*h��-)^�'�q���s�0��Dj��fp2�Z�E���ڵ��lB�2=��[�=��5,
"!l)���Q ���#�F�xT���lG�ԍ��)�$��Bי����+a"��@*dC7<g��e��w
ܬRn�Y��s�%kA9De�=*Dkx��n魹q�:;���A���+�1�Օ��[�T{^�%!?�RU-�Vn�"`K}ȟ%՟�����ZB8	�kEH��ă��,Z�SĪ�8=x��ƽ�
�(���D����_����I��q��:&@ģ2�u�G]amy�b�������A��ۥ��%�\7'L�R}�~iX2�Յ��� ��+PL�!�K3�\�G�f�鉽�>�����n�?XB�-$���+H{��ײ�r<��5�~���z׶���X��Z�fA��MS1 D 'b*�",��u��ޗc^���r�KI�' 2�[�hO��x�-���ջ)u�i�?~�U��t��"1j/r���7�vMdxu�JѾ��3��B'r's��Q�,"���meY�q�Xl��Ĩܳm�v��/�RCI�����nf=T<ᓻ��c�C�(8e�A��ཕ&鯅*UcO4Mv;���,"�"s�s�"�8}��r���nr����1)	����Qï���C◒�+3� l���۰#��ù��T�g�B�_�����#����">������(�`�Aꙁ�G�+(�g�}�j�P�M5oߎ��1<Ա��hZ��Ѯx�H�0S�|1z�m���ڴ��' ZZ��ZsHZ�5���^*�<�,ŧw��d�-w���ŧ�a{�� j���������KYe:�����$"ތ8#��絗�y����ǉ�P(g0�{�[�6����ܷ��SoN5��Z)�#�8Id97�W+@��男�;�
�|E5�f*aK��v��bävH�85P�x����tc��#�w�J��끈eA�deIj�� L9fL=IX�۟��g ^�����ۡ���ο�'�w�e�
 _Ig���Ho����g���X��(����������Xt����.���GT\L��l-ބE'��<�T�hWO��r��]	7�G��KWz�dya��Ўc����U� S�W�]���@�*@�c��r#{|~���q:.��(@PmC�{B~!��O�Vb]��,���|��{�	p0�HЃߣ�"��������1�f>�Ѕ|��hp�][-�P�Ū��>0��W�O2��o?��f�L��?������I������3nl��O>4ƙOb+vX<���_�{���ҖKu�����$z}�G�}h����@O42��_�1�iȯ9ň�Z×��V["�
~?�O�x�9�v�7��GQ̈�lh�|��3������M\uV�>&�������s���U������I�DN��y9�=@c��ֽ�%�)hl(��3���=MK�7��#�c�gT>��X�pzT���k��>�s���>��`}�*���tn�[}I5H�0H~����p�T|�%20�UY��j��Jx]y�ARO�.�i���k@vU�/���0���A"�=��`�yWs�S����K�1=�xt�%z��[��%�e�֌<�ڋ�LP)�`���?�X4p��w��	�:7c�?�C� �G����O��Y�49��
ǝc�y8'�x括f2�������⮊z5�(J%3�v	B8��d���%���@4����g��9R@�䗛��!�r�*q��=ܝ?|B,����to�{�D�{�$P�3ub�K�����o��m��y��L+��$��0v��bТ0��J
[שN��EQ,7!��i���rr7�G?�?����+HrmɃ~-�J`{��U}�:O_�B��6�P��ZoW�\��,��oG���E�� �Wč�0!�\oM!����^h�)#f����B��F�o4wr��_�_l�%��Ɂg����(į�t/�WU�8�~+��'(`hȈ�yᤚG����������L�H;���o㮞S��IĠ�p���J��U�k	;�e����ָ����vŚ�����C�Es1��(a�!bc��0��?�;ki�Fdyj����i!����u���#�\u��֬� l�p������6�H��+��_L�Z��N2���Q��^���\O�_;թ\�֎��FtRqN1U��HS�L�F�����_��jP?��{'�g �R"Km�VM���(���` ����ԇݦ�
��*uX����z�{��p����x��T�Gb����.� ��^�2)lE���G���ϼ�ks�3a�z]�.������i�g��i��g�8�Z�e!F�#��ⲷL�
w:��W�
�r�3��A��sL�d��}�l�#��`'�rU�Q������������O��S8���e����⌚J�����	Y�i3/N�jHtC���rOP����.Fַi�%SK�.��]�]��~6����!$GI�"j��|���	�XN3q��i5��q�1�@�|��	�#^�����T`����D0ѡ.͹Ɠ|���s�ß��)��@�u6F�ζX��pVF���0kf���(T=>]G����1v۟/ʌz�a�j�[s@8��㰯H~1���=M�92S���Tf�W+�m�i�/�q�Y]��/�9>O2Bf�tj���+E*ֿY�.�B�)�����7�ݫTt�̩c�V��v݊��SB}ķ�T���]��[�)gPi�D�䤲�����E��3�˩�Q)͏hSZ��+�|.�6�5��&���&��X�9pg7EP�O=;��R�ns�w�Lܺ�,t	̃���h7��T���a@�`T���ђ�y����.���C�O'�z���M����@_ɘ4�\�o��z؈'4��C�����3<��s��H�3���Z�e*f��_P0�A�J�%�~��6�%{�����n����|����z)��蹽����0��3��H�}��e~���]�{�8D �ǆõ)5PБ$��fWǅ��0%��B�o�8���L�6��
7؝�o�OV�tr������ύ-�� Z��6Ǡ,�3q`ʜB<�%�b����fRF������C�↵ z��x$LNyM
�3v�[b�> �����!GGk���Q���#s�'�A=��TA�T1=�X�D��^w�*_|�&����ض׵��`��%�gWq�W�t���*NS�n�����I-H*B�� ���`ʮ�Nhd��r߰�b��F�ޢ�<X`y��n�������=�K�=������:��/��~�yx����ch����dQ�)E�ũ�;�� ?�� �f�,ܩ��.B
��Z2�$�J��"���!�(-c�"�����a]/�+���Z�aG�5��߬�Pm�!L�tt���
�q/���469`�}#��=���c���z����ƶ+�L��YM$X��j���0��_���r��Ѹ'�C�/R��%��k��:��j� ���s��D�v�`?:�=�9�q���nD�5lPXH����jJ��e1-�(��/����E��2��|�����=ML]A�rÐ׺�=�%�3#d�w6�N�/���,� KZk�6���K�I��&BGf�x^b�4@F7kT��栘	�ʴU�u1���6ߧ%0u R��V�pM�_JJ�)��3;x�X�{.r�̬�����Öt�o1J-���co��m���AYvph��G	���n�m��m�@�,U�����ÿg���!�r�LY����oR��s�4w�擋f.��i���u����ZOu�4�`z�3�ur���ȕ=j�������P슂���Oe�՘t
����B��i�YvHzZ|d����۷�{tW7�b�r�v�ػu�V��zC���i���ֈ���B�ccZ\����HL5�}4���.
���'�=�5�Y�ȴ���R2�8�ݦ��R/���Kx�&�
A�J�$�e��6��OF4��J+�]h2����d�֨+J>��a���a�ѥ���s|ܱ�=���g�����.i��
��d�����\j[(�4���/J!�.�i�i��LW�t2�I���)��-1�#���)�S�f����g3���Ù%xN�P,��P���<��_�0*g�MT������t!E�A@��#ۏ[�L�;����|���.[�]�������̈e���s��"+�N���j��x���hO�<>o��M���j  ��	�E�$Z�Ј�$5�1�0��^w�6mh>
Q]����5	�DA��1�tW�/�~���c'V��h��9�~PT��ClE$V��i)N2*��=�a��N�<����}+�#�^�2|�#p`#Mf�a�|��T;�Y��O�4S*�W}�ğX�j�v��|�u�:�e��.�ϔ
#tB/U�Z���RM�*0ČYu��s�0
y�1f{<2�w)�@T$�~j�T��(���K��&ɽ�y��*�Rl'���9^ .Yu�8�uW���[NI�G��B�J�~}�>��f��D��o���H2	aE�(j�k��n�MR| 6$�	�䭻�f{�U�g�<Ƕ.Su�d��U��/�F3��n��������}�VA}$Y&�W�vZ����J��H�lP*�i'n�w�h\O�=݃��_��*�}΂;�o����i�x�c
��l��M'��ѱ�;qXe�+��.���Q��"=���AZ��g!!<X�+��%P2�����V˭�A�Ð���!�r-�5���|� ������ ��m�&�H>Jy��A���@ڭ'�\oD��@�/���PZ,�KVL��.|��8����KA)�MЩ��KlC�$���O�2���5�@��hl�8���"�XBF]�5����=�zb�j�F�O�� 3M�V�������,�8��ae���Z��ȿ����*�Jë� k�jR;<~�,�X��
bt#�D��K�nq?g;9��T�����bM`���eܫ������ue`Gwܬ��D����I�ѕ�`f#��uD�? �r	�I��}���-/ ��\�gT��?�R�$]���&J��^,��(�U2�XRin��>���W�J�3����d������]�F,��D@ ���5c\*\���UB/;��ǂ��j�>�,EU�̯�j_����q9	h�-�6ņ�x}E�P`Yk;��
��0��Pܱ+��ڢ[��Y���o�9��B+�r�hqs��J��0���-��0���ujɫj;���;��g�n��:Q��윉�qo���"�8���:j�u��I:,I
V� XO�_�Ξ�����?���ubg�s���ndxk��q�ǩ�@�Y0;��5xT�Q�+	�V���a�rR��ߜ��\G<犼%�+Nacխ�!-�ϥ�i��k�s��.��>#��� �~P� ��u���ރ�mh�5�J��n�H�<d�F�[b���xͺ��Q4� /y���^���C�R)u��%����Z���A�y�5�U��ŠΟ���x}�����nu��[jPY���v��A�=?c ��Utb��E�Qm,�9:���j��-t�Ϣ_V�(�Ů�@l������]_��%vš�h+�'�wY��f���ߎ��������%j�:.i��|~�%���Z��J@�R
5�
[cͨ
q�8��A�>#gl��TW� �tïO�=U��ބ�வ"�iv�s���s�Ҥ�����-~Nhg�u��LL˨3� w� �\(���ˊmݟ�V���&ĥ���I����V5�F0h�OoXX�\;��1@���]�p��AԂ��GG ��/���DY�D	��H*E�b����P~I��� ��DWG�7o���|笲��rl%8����Tcv5�B}SD4��<ù>Eϲ��g�U���5�h>��Z�^*U����U�%e�
V����
����O��r7���sdg��������L��
$�G���M|a{�\����S;�]�];J�^���6 �f�L���|,R]|Й�ڮ�����ƙ����A+�!T}��0�L�����˘⓯��#y�$�-��^�>ͫ���c;S\����!3r�^�_<���8�h~�[�!ps��ض��8��Kܦ�%_A��ӓsE�ȘA �<+��<���|�u$����	�	f\L�a����8�|贗m���>��k��� �NGC�]+e\z���9lۑ�{�ǳ�B�6d�����z�C;�	����������'��+�G9�!�-Ạh����uV���s��Z`����o�������,
n{��\����:�X�۾���{TT0CN1ۀ%_ss60MG�pU�@�r�p='��_��pN��a$&YjQ�U{���in֓�mysZ�c�"Q�EyCN�xw�����,~�IY[��.	�ѽ���U���:�(ٰ.��E��I0�+����
��G�n����^��^G�{\�XAK6Βw��֓�?|ə�?����ؚ�2�q�`�� �<2�v�G6y͗�'����A}w=��	��#؍~.�G3KGFlsz��3׮�!xV����B�(#ϗ �qWM�2�e6S� A���ߓ;^H��^W�˂��q����50ՙ*&�����ߊ�rIʼ��Yt��d���(��z���[��+#�^w��b���Z5����Q�0!5BRxQj=8r!�< R��!Q��5�Ϣ��J�,�����w�K���LR��5K��Ʈ��SlHJ�}j(�&�$RE;o]�h'Q�ǫ��ɤTyo�ݿ�#_�����(�j���7v�[]-��2bCxp�DN�����EC��U�9�t���h=���d�o�WŎy���mg��a9��]c�Ge��x���uɱ�`+���J<R5���V����N�ikL��I}#/fmD��ZgE�U�u���E����(Z��a1�^#.9���Uu��f�5/�d1�H2"�Ȳ)�p�Ǝ��p�	��^��>ʍ�rPjxP��R�l�4UG�9Y��`�t�݁�pV��|�7P������c�G�%Gn�Nh09՗�<�Me���G��	N��,'B�`UP̍ө�~�S�*Ɏ�v����֩!�Z_��-
�HHR�)@Fw����d�낙�?�
��hT�,b���#�bU�/Ho�N��x_�G6�v��~��ab��3~��Wd$/���v�m���*7�V�����Y��9����7�o��a�G��j�|EXt��Z����*��3�#G��vn�00�3��z�k)9�)��	�<1������DL)��U Z�8���9�#K3wfYS+�6K��C�X�oz)6�^���o�F���}�= �;�	��B$U t�	=R��Yt��-j9Xclf��zu����\�՞�]r���i횛�sy~���F�y]�CfG�؍��~�cj�qc���q����?ʀ��54It�N�L� ɖ��m��>����٧�+��_ў��~�w�z�KvC������ӵMn(�<1��8®����]��'����H5�gV%�nyʪ�_�߅O�6��z���0q��,��u�Z��͢���s+VU��{|r��Ȏ����7 ��s����L�	�NP�26�y3�
