��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s�����׮��3�9 l�ubHe�ዌ�K�Ey��3X�J�Vϗ��1�ð��(5��[D���v�C��"B�ݶ�[	�c����}���I(q8[d�UB�@+1к�VBy�%7
`�5��!�
�W��ov�@d"�➮K�%����
�n�x����\��� �qe|	7wQ���:Ddt�5�)��m�BA�O��m��*̹;�:�^�z�l>Ta?coP��O���}��mLU�D#�s\v��v�R�J��8�L��7o�P�9�u����t�ϟ���HQ���6В>e\W���9<h>)�$��D!�C8��H�䮨���w	�H���99�.9���-�tR��;.U�=�xg4�]��#�->{4�0�{{�=�M5�p��ðݚ��}_�� A�Y�`�e��*���g�����hϯsg-��u���0�R��Fo��za&����G�j}]����LF�������

��3H��ZG��$qD-te�_���4�����^(I/V�Ó���иm��#���xۑ�δ=��xq#��u7�T�%DY`|?�=��*�O��_��u��;��!`�^?�0K0U��Rg�.�<���ER�}H��{mcrlt���6�j�g� 5;/�T���M�5LA�Lh1��݉��.�ກ�5��g%�eQ���Lr�m�ᮂ7^8��ђ���A�*<A�.��ZpC�2�R��/g<�L��=�"R�?/[���<�`r��`�$����C'��T�C �L�j���C�|�#G������tW��55�U���0���Q�"��#C�V���,����7\���4{�ú<;�T����1�3'C���+li_�:���0�����y[ˍ���S��q��*9�X�ޖ2��X�ǁ�E?y�핣���]�)%����*ti�sN�b4N�g��j��~��������R�婑V���� �vC��a{!����:�
���1r����s��W��b/����6E�bU�����P��v��� �<�^'R�^�^H�d�qg�u�*�0n�I�νP��� ����:�{�ơ���g�����̫�����5������A�"�]�њ���<��H^͑]P���(�iM���c�l��W�J!�����b�>�-�)����X����O&�<%���Z���K�����00*�6�NY��Lw_v����P���3!ѡ%��S���7����ǽ��j��V|��7Ո�0���v�=�/��.ebxe�Fw�R��,��W�T�4�e��d��EI�=��Q�c������F?|��%$t�d0����:�Q��ù�0%�\�;�/�O��j<�W�����%��p���Q��/��O�q���f<�r��Ea�9�ު ,~�Q03�T��Ox�dԈ�CM|�Cy�	?}l`c��fPwN�s�3Jj@h!�}�j1̂�վk�$m����D��F�����h�@�s/Y�t��dĺ�����o�-�"�y�EYʾ�����p8�k#����V�s0�D<L��<\���s�#�U�u�����Λ��F���ʳ'��s�F�xG�uї��B��(d�	���  �<�� ��hȹS�w5��=5�Kz�7�|�i��Ԝ`���|�W���&_(��ޗ��,�W{�!�ҍ�D:���-!Y�#R4� �yZ^cwÖ������]��0\��W���cHQZtO��s���q,Ы�03%n�6�s1��D`[ q��|/%�<��?��Ĥ�S�:ac�a�t?~�T����!
�/�1W���z�`h��rAr(R��6'���%Y��'�b��O�pG���0Q���~�З0<�� �3*G ́����?� � E]�T�z���ۧ]��?j�H�h����qH�+�8"�;�r�(������8����DKt]�4Z�v��l6\ZI'�v��޶�.�!��� Noh��K�i"���y3�ᮛT�=�G����1�%G��	ǒ���Y���a����+���>��9t�pi�15@�!����Yn]�0���eMTD������,T�׬����D���4�Ho"D��ud��<�,;���԰��
,|��iݕZ�ܒ��+�0_N�SQC�y~��c�dN��SR��*N��ʐ�(�
�f�τ^j�K�b�}�|�-<c��=._����o�~wS:���2�������Z)��~��d����nqb��V��d�֜n�0�f�7�[)���o"�,A�<^R��ެcH��3�&��H���̏�N�p�,j2�Sh4~P�/���������L�P�\h�_;S�&�K}���}]�����"�S��U`�}���
���n�N�ה|��������4�:��Z�[H��/eRST<�M��R��/��e��GE�t"���9��^f��'"SZ�g�w�o�aj8�ԋ�d�8o��T+�7��=!��o���������<3� �a�H��&B����a��e��#e2�R��co�� ��Đ���?��I}i|NW�%)���nY�kh�8ыӺ��Bn�ɓfcT��]���@�G��qQ�Y*�������R-*�"�&�Ќ��6N��t���I&�k=x<�C��9�&�o��']��ڹ�-��Jbd5��0�fVs_�Z�µ���Y+$�O	9�?���FIZ���4X�kg��K[.��)���w�����pMw�!�y�z�0	,*vG��<��&X���E�i��Omo	vpHm�xQ�L�Pͭ^Ȥ3�b%����@�;ٿn��P�cA��.�6���ٶe)�o�a\�`�V��Ƥ	�Z���槰���ßȇ`�I(j[�|���!ݢ�p�
�kwL�V�E�B*D��Ǒd	b���"
��I���x#��$6����If?�
�/��6�;L�E_[��*�6���p�ڋ<����}���	���9k�a�E��zH������'����}�����Z� :S��R?�>Y�v6�Rx�ٯ�= �{C�q�2��f���K2
,�`u��ԡ)�H�1)�L	,����:���t����A��f�~*��p��'يK�$�,v���I�U^�\�E����	"�f��=vL����8�Q�|�IɄk�9�c-ͅ�>PCR��=�Rt���ҳV��c	!ڠɅ���2]f������*�Zp	 �����~2��@� WqE}�]���\��� �6lI�K��H`ؔ:!�.l�z��Ad\F�{�-�t$��\�Y��;+�7O.>��x�XP��\HC��6˺� ��S�9p��h��_�B΀��m1b,%����u��w!����B�jC@��:����^��6W�]�2A���tU��q_�X?I�ɥ�O͡�BStf���4:� "|�J�Yk�$xi��ξ?�u|��������M��H���B'��̒ ����h8��"�������y+,o�CT$�]ӑA�. ���G��b@��:\��y0-���A��kH�,Y'�{2п���B%6�ŕ����P��_��۪fR��g�����J�	�m12J��S͑�*@��O����@@�9u�o��dC��#�$m�K�����*����!Yp�35t�ೂ'�	��UK�KܢK��s�S����;k~W{�3�)��9�$��4�-���;݁��#د�H�1A7�m���<�L��C��$���"A�jg�5������?����aS�l�ZD�[�Wm���Ѯ8���+�� �W����FYOZ�k��R�Ypz�j '�5���3����058�|��KB	�U)/�G�>sdv��f��K $��ɵ�Fiѷ.pK�(�eQ�h����5y�w������h̚S���!�m�@�=�(}�M�Ŏ��vvy�Yo�o���.p�ڌ�
3�/�������&2��?�ׇ��L��n���V�>w�Ŏe0��9�V�	0iG�q�넳�B^�	�X5����6Q�G/S�_�I��\;D������[[�a\�{C�o&=O��@[���z_�Df)��Ҵ���Z��ڞOH�z��CA8b<��ơ� ��,4�עT�Zj-�,�����%�2��#u�<���l;�9�h;�u��,�ɬ���c����G�?��'���y�/�c�>���p(��2��ɡB7��� R�'��R`G^g�@�Q`pl^�v8���m��W�I��/ `��BV��0��75���]z�[����������ظy.��L箜4�M"h���Z��!�T���9A��̎|���Fzu�/�aM�d9�GE�X'����2YcN?�'ϓ������z�u�~�	��4��ч�$�������i���}���$��C��I_�-^'i�nf���⥡:.�8E,]�s�W�/$�v��y�-�RS��%p�<����V�p	|�L�7+,A��ҏT�ס� �Vlѫ��yy�<��_�j�܂��-��m圂��=e\�ş�:؈+z��sݴ��׮��sB�+���)H�7�`�[vJ��M�)8(/а��D>�&κ�XȌ ��&�rɈ���μ`�m8�,+�����rT�.ټ�T�b2G}zk5�ѐ,pa������U$sU�=�}#Ja[���ٚ=�q�ƙ��&��afP'����s`��{�4�&W�OW���]9�;?>��l
" u�#i��A81^rܹ��j�+/���T���ș���.,剴����b�C-���<������\��Tz�1�Ai�!W>�F�:|i�3����u9��t0���0�fH��r놄��24��D�L�xw��f�z9G���zIL�����Ѱ�bO����M�I�����`�[�.��t�+4,��m��������վP�_D� ��E]z�(yi�:q�/Q��`��K0��� 7l������\Ň�����X`�4��ü�����[M:�n�&��y��V*v�[�])�U44�jx��2�	:�w(%s���?XXl��$n;}H鹭�n����=��?��;�r �� ����+�"gd/b�8��.���o�>7�G�gK�����X |xc���;�GV�Q�7�D��{Y��a��=��)ꋬ�EJcT����_�B��zehg�W7�j�3�l������ɡ��g4����LM�9��%L[;�̦��fH.<���}��{��{hg��x�Y�ҰD���/y���0ڰB��Y[��EXSPz��V��sdF�x$Zw}�d�oS�[L0}2�_��Z�y��8��[�);�~�bċ		�`�3y�<x"DW��Cԙ�{Т{i5��=�ߴ Ÿ�P�zx��P
�Xj�֕Ɨ�/v���WSE`,(;��J���	4�/iS�M�E�Z��5!�K{����oI��;K~�U��"n���J#�
�:ˆ@ w�K��vu�B�'@X�c����4�4�R~��q�R�`Km8ï����F�&�Y�}��3�P�_Ml��OGi�����/c��2F��4��WYΣ�I���6KCkvO1�����J�PVg��\�:k<�
� v5k���-��^�%T(��䖅ʧ��;x����d�ϒ�
:�~R���ɆQ�eN�P�DA��{�e�+|p[���c�x��b��z`Ib�q% �����UH�X�Ͷs�:#
,����S9�4gs;�9e��fT@�i{WͿ#���.��t]綨�Te�Q�7�Z��w+��4�S����v��u����f�5�K���Gj2o��^��(���ђ�,ٓD:����_)��Bdr;Co�/V�@�q����(l1m��V�= C�wd�}���S"f�U;8��� P_��gD��H�Z��0$x5��U���W*+�$ԯ�	��� ��zg؄����!BǨ�:�[��6th�i{$� p����"P5���&c���V� ���Cs�����.}���U�&טZ�ަXp&&��t;KN�x���U��
�p5��-���`�ASk8�;S�n~�ذp���5����I/�0��"x�o;B&g���A��}��t;w�K���CYGs5rO>��[;�I�3�U������iʬ�b��kt������}?2{=L������;V�=��Yù-����"I{	o�ڑ�ZX®g�{{,�HM�X"35�c��Z��؛������'����x;W��ʨ����~$�p�����-������c�w�����r�����H�6�楜;V��g��k/}+�Ëћ��݊�*-�������|R�:�3w�ޟ��oE[JZ3��XagPÎ[��{?�7�~
?�]�F�@��u�˫ex��-�,ys��["�	x-V�꟩����s�K[�RȀi�?��d�|����
n�R�`B��p���xʬX�*�&��?�n;�n����2m:�Bw���8�H��1.�i�cX(e�D=l��#}[U��9i���p�W��\�4
��H��蓨n�Q��lXJ��P&"4{W͏|����PJxѥ�2�	�eԏS@$�b��ʂ����Ȏ������
�䇭��qY�5~oz�Vik�r�؍8ɿ�J=T�� �!�XY�P��=��|t��\:��L��gEأ��������b�L��%^4>S@a_���ԁ	Y���vh���� ./��G���%t�ұ�)~VTG�7C^D5e��Q:W�H��8p�5 ��2�S9l�[��	�
��=Q���5C�S#��G��F�]r\�^��{
f�|��f&A���p1��@V%�;�~)β��;����dT�m����}T
�BI@:6M��诗L|9��7+�zP�9XB璆9FH��S�y���m���MC�|�o���}zi7+hI��[Z���Q� j�,u�����:~B�?"n�<sԮ��t����G]L^QL�l~zqQ�%�%o��p����=���|8 ��P��m��s��h�5��-*��)3��*=oƟ�m��g���Vqٱbjvv��Y+�������!����I8�'S�aN9�ev��ݫ�*iƵ3��O�#`��{�~"'�IK�HZ��Wr����x��|��-��9�N~��!T�w���ȧ5vC�
5�:��k��&*�yr�6�:���F�	C�ၮW��c4y*)_(\��e��N���}}�7V83˽	�"���v<�?�=���e`ǯ���r���V�P�J:���M�ж\�#�X���r�X�̞�8�yI1��v�v"�f�yV�_��W�-���/��o���]�3��,���/V�H����`x�n� j��R9���jh�CA�# o��`쯊Ө�E6����MК%r!'�([M�"�g���1��������)��:-�d����5,}|��ހ�l�,uE��Y\�%��3�T�8������06)���w@�D���8_�8wc�^������pG-�W�����ݯ����)z�_���QT�=�&�j�5H��"`2��(���}����'�'�չ%Xz?�^B��S���r2?�"gH�
Y�(�Gv��aR�=Ds2�Dݵ�g�'~RV2,���b"�[���c����1��U7�\�`:�U�~�'WB�;~��)�W�ѳ��tB�����(3)�^��6l�X��n�7C���N��:<H��(��O������i�s�\<����{�n˛6x��P6]U�g�1��6�Y�3k+t�L���� 6�$�`=�_e(>a����R��?��ށ>�����Z��(@R��������"���C_X�M���q`��@:����l|W���$�{�sg����i���F�Z*��̙_�U��q��)[$s����	���OV���_�W�Z.
��v��_�s/3���?������=(��e���Ndd�pj��D�]by3�����<�ŧH(�̗@�Rh��vuM1(���p�P�Mza�L;��f=E-��X���a�Ţ�{X�ɷI������o�����k�^��׺{j1Ƹ���&�z����i�_�����Чl!���t��|��؟�z��e�9M_B�P��BE&�tn�����=��l����]Ec[���n�$R�YP�X��I�i��^1�i����������p���� .�{�A�v�6����Q�t�݋��:��5'pZ���m�����% �c�A8Q��_0�+%�6��;*���T�߉k�B��n�i�����$��u� Ӄj+�9��^��S�\-�1�̻SC}t^�i����pB�2��,m��D
����ˆ�*���L8�.�P�a�Ʊm`bR&��7t1b�3_����ߖ�����Z�	��i�EH! ���F	K/��
QV�)�]J��Ƞ=��m��V�а?���S��uz�՘)��#r��	���N�S5T�1O9���"�ܭY�X�
-���x�h�\�[c ����jVot@����; C=�h�M�U/j�Ѫ��230���7��j���o⓮.���}�ǖ7w��*����M7k��;��sI�+4�xe����+-V��k�潨:�Jʝ��TT4 �Ǆ�N6v�'ަ|����-���CY�E�t��Ҝ���bv���3�:4�O�\��Ȼ>����_�;|c_��8ZX���	a)ƚIj�T��C>-6Q9^9�r7%Q&�f�X��fU��&#��w)���X�ڭ�T�������Ã�7���J��2v�E�����v��((�5����������� bs>�~�sPe�
�O�F�iP ��Py�]�����Y��e��Pv��4�)�5��̴mx,D�*�wq��>�q�۴$ǧ�!VGN��:�Ha9���b�G��q|Y��+��<�l��C	.�,w��n��c.ʵ����W�	.x88sLx�Rln|�q��7��*`��u�i�ZD����%�A�q�x�{ߒ���t�3G�.�BN�����'=�D�V���#��D,�O'^n��˥��Ζt!�i7f�~<ZT��f�Bǳ21����܅��1��g9����ہx\U~�Ͷ�&���NX^��'�Gʔ%�7�t�0Srz/��ahH���i�6���m��jޝ�+��:�R�{��F�|�5:�}�<����%�]��F��"%�u�5
M� �zyw�ϓh�VLc���+�B� J���{HHК� �j�kJZ^&�/�7�n��(Pd�;1�٘P^?k���G(�����@9�[M�m۽��\l�z"|��-��96�S����+����%j�Rs�<�Ho�cL@�w��Y��cl�J��hۤ���4�?
-��0.������"i��r�qB6�L�
�5D�<=��g��Л�f-�w�ׁv�^IImDz�	v����!�ւ-n���a��@�L���*����qD}d7ch�̝����uNz�.��~�AE%p#1��.M�h>P�԰ʼW�|13!�7��*u�l���"�.%~a�������}l8~�� ������8���r�G4������mO��֙x���Qkh����*>�{��(ٺ��&G�|D�k�T�q��kZ7hT��I��C)vt����A`��غ�T}���5��J�*�m��S����)�0�"-xdԣ��m0�o�Y,�W���I�'�+��7-����5_=�6|	��Pt'��x1=늼N,��1�[�֙*�Of�>BC>*�X��RAQ2"%#�@Y�Љ�)3�#�Q�ކ\�Z?oy �7��=�&u�!�We�6"��K��Y�Y�R)���B�N���j�G<�˙y�_�� ���*
l��+*�����"��U�ܠ�H�*fI�6�ƖWl^��j�[|���y�5�<_�}�Ȩ�n����5����e@f���=� $��#��A[>�z�&m�-�֨�瀦�Y��.��%���JT#�eWfNv�)nv�<_�DD!/�F���N��&t�t[��C��am Y⬧����0�~38玳bI	�J�����EC���U�#ήTX I��
W��g�tD(��>O�9���;��ܓ��0S��O��]P@� r	DC�e��<x�29Ɔңzw�>1~�C$B=��qxfz����~��Mj�Yy�tK�?�>�Ow%�̡X�Q��ٜ Z�DN9��^2�	�:w�P��ɪ8�fp�V:W�9��H�8��6����P�E�}Ѕ-0��8�U����܂��Hex%y�:R"��&���P�0*|>���f@�����2�����!��GrMfS�6�js(5�+����F�5��Uȡ����e�"Es�ctK���߷���!�s������#���U{fO�ár�$�
���i:)h�`N�U:U<�^@S�jmF.�6@��vW�l���#�u���X
�8�3��.�W�[ ?���`�����9�斬VT��)�ȫ�� c��X�2,N�#�J�-�nq��G��Fm#�9~n/��I��v��j��쑘�0�A���;[x�z<�5���..���*��ᓭ���*>��gY<�|�ac
D�G�B�L�i��h�S��{/g�*3��a_k���rO@��'ɂ�G�)
����\���h���T4��m��3xO>%�h���iG�CA���B6V�1i�O1��M��גV�^V�q��3��;`�x���vA���'o���R����h2�b֝��Xl��!��'s6�T�;����B���Ȫ4��~@:b۸�i����H^ ��0(��]Oul���t�Y�H��庑�O�,�>𭂵��aԋ<����/�soy�e�Ė"��
�R�+�`+���K�A7��	��j�g�1镪��ج
����+{W�!%��\F���Θ�[&��Y^��S����\����G��F6p&��$���)0�q��!5 ��j
�C�<7�^+>�#
/���s�L�n�>n�>ߵ�����^�1}
ye��_xG���^2�JQ� <���0䥔^3�1�1:���. +?�:��q����k�X�ԣi�ݳ�L�>��AH�M���%4��<T@w�L��J���D��z�u\Q��&�r�x���	bgF>��%eft�bg~Z)�2�b��o@��j��U�<]gW�j���v�.5-s�&v*{�Tu0�
d:f��<�f5�M��Ȯ2Wm.-Z4����=��׌�o}�̙g�2ah���{:u0M�|���(,�ǂ�9�˟C@&HWi�v�j{��L[��YY��иᦼh�P�A��bx�h�39lrc��������S�u^������TV獈��S�ˑ�����fMũ�\��XU3h��$���a�ڝr-\����Ԯ����ʹK1��$A9����$�8Ë�!�5[�D\5�Y�/_����V��SIG>im��va�=ş�q圄��� ���j���t.�KrW?HX� ��Zy�*��j�0�J9�nγ⠠���C2:B�6CC��@=N}�:@>p��8^��Ꞌ�p��&�7����/"��Z���[]�Q�ʶ���o�
_�����&/= �گS&ڸ��Ë��l �D!#���H�!�0X=���.qI�t�s���f�|M�.YP�.�C�6
ح�љJK�FvOX��H����^Mi��g�|��"�m��z�x,��s<���<�)�W���V2$�AL2贶��������\!���Y`Z�L�ݼWm�5yn���p;+z�����{Ǭ=3�v���76Q��n3$�
�b$&56�@�-���1ar�+�$KJa��;��MS�M^$O��a~ȣ#Nw�~���Լ+s�p�B\�v�C?�Lq���[t�w���gԃ�=z^��У���`����ӴM'.� �1ɢz�����h�v��Cz�����ɠ<TRƊ:��t�5�`�gLO�ra����	Ǝ>�����A�̔,<�.��ȌWݖD��$|��3�t�_\}���^�E��:�,]X��.o����7��<�H�ѡ
���VFf9͡���j3czk$�;��<����{mYU_���3���*��7����a� �|B��iKX�S����Dx�y�2���F1�6|�Ӛ�2'��Y�,�b���$�P֝�W(#�:�����W<���J�pÎ��:�(˔.�[����Owf��m�վ�\ �G����I��*���({�_	�����^�3�1K����A����r�A��#�~m=���� d-A��]��3�1���d� y�U�^��`d��`���� Uz�Y1~�� "�l�q<+��6*���e�q\�D�Pw�I�,�^]g�s�'�7��Ji􁛉��������5>�.jX��zV�H�� L��*9j�PJ~(z�~�޼�Nۂ��K��	�]Op����[���vih�2d�/V�o�q�f�v�x����"e����~)��n����`���_F�#������x?c0|��P+^��5<T�	���2����u�g��{�!X�O+�G�ݿ�!�˱d�xZp:=b]{�U��YX�0��,TR����2��S,Dc�ҏ7K����Y����W��˺�^�ll�I��gW��j� ޯ]��)��Z�xCʰ��zɭE��bR��8ڬ�:�|����۶�}"$��f]��o�����S�9@rĈ����y]5x��ײK�PIݐ4�����l�����945/b�疍�7n2�JZ:��Y�mB�N��;x�v�z����-u���9�Oc^B�R��˞���+�l��,����o�d膯��й���Os?��.�K�I�}Δ����@N)H�\j��a�k����H���s��-C�λ�ԳF�x�?�n�wF�YK��*+�W��(@�\��B/G��l�ZE@߶f���d����>��E�Tй|S���4���rw��],AǈF)����`��>�8���-���<"�KM�{�k����j�w�ĿE�[59����5���1��t1@���-�˵Tj����V\�Kj��s�wgF�ǯ����� e5=u��jd�!R�-�]�C ��:噠֖2�F����F�$z��'�y�s�\�3����VY3q;�n ��������p��~m�~�$sZO�-�����d�f��R�!�ZˁchkW��^��^��0O/��=wjp�ͅ�>���:������U`@�C�0J�E&�H��9��V9��㊙-c���^��|��h����d��[�/zO�W-�_ft$�aV�JǒZ���p�U�4JC�
E��bN��|SEٱ���0E�	��"��C��g7�F/����Ȓ��@F��,�)�Op<��%A�g�L3��c��K$j���yt	*������lԶ���,�3`G9p���ɋ<��Z^���uI��H.Ž���x���b�lA�gM�nR�1J���_����n���O'u�(��u���;q����rf)iZ�Pc�̹B~��3��<xT�`ljA�z�:���M�N����,�"�%a�E�Uxa���0Tl��]��ȓ��Z�NWG(����3�J>p�G�ɟ^�����u^�y$1S���P���!L�m���k�@��Ș)��� 5����<j�.���"��r)*�Q�4Y�~�t���8~ �>�çgY� ��`,�N��伃E��.!;��g�V��K����R6Ī,�$��4��|�	�#i�.56�I�ihGt/��$w�
��5i&"���	ø�L�JoI��A�G.�1�B�i��t�W� s0�W#�ﬞǘx/f<� ��&@J����4����Q
�딖��tV	i�S��e�F�(Q2KA�\��.@������&�	�bxD���u3�0
ȹ��ۮ�Ă 1�ľ!;�8�=PQ����n���^K+�����*S���Oz�J:Ǜ�����ͷ�cV�%���D���^�Q9�s�#�j�H����Tl��W衩0�y�C?5���|���y+AcQ?AuYeoH.�tz{�k�:����6�w�T���H OA�c��f�o�8b�<C򢁙mVTΣ�k��A@m�%4�Zk�o�|�Ҭ�~��bE��q�
��&7�m��؏<x<��]P�cם����#�>ib��֍�K˴����i�?�#-ƞ��	�BM���3�j��0�MI��>��5pG��eQ�m��\�5��n� ����z�v��Ӳv�7���jK�"��(�O�xn ��M2�7��~�&���!��3����©hF���Yɥ��z�*Y���^ϡ�r��
l���-1�n��J�����?y�.�$[z�Wn5�ΝY@IH�ʬ��@"j�ӍM����<N~ �<3�Dh�>��|/m���<e�<N��O��C�Ȗ��P��#j�&� 2��&e�f�*(ܤE�b�h�R`��0�O6|`%� �˹CpS<ؘn��
	Q������Y+���z�̋}�Ƣ
�[��.��:�i7����b��E2I�����@��>^7�D�i��*y�bS:x����߁���y�P�e�f5�Y���q��N)��'n��5{���V���x~w)�[/��oH��zM�m���md�Er�{��;��2۱p&��M:��s�Hp�W�䵝�9���P����+/�Б;+;�l��G� ���m��m5���K}(�lPfL&��WH��7�8�}�+Ok��7���h�T�����3��AO�g����v
3��n.y��ۤVENנl�"�s�
'Z�"0�`��m�x�@ќ�E��xJ��W���к��%��7\����'<^��5B�#�2��Ca�^W�}����3r.��1���v:E�r�O�[6�:uR/4���/#�����s����)w�So�(�Z�k�=jdj���A6����❐�а���\��� �,��Ɯl���B�ZL������c:'�|>��9�d8{i��f6ǥ��J{qs���薖ӽS2�8�r����?�^(̼����ꟳ�zHk(6w���]a����"�i�Fg��R;s����X�����+΁�bb7>�h��/5�wx����oY�q�2�_��e�>O`�O�<��%`xmk�u�5���+���5�%3/܋�+�k s��#�T���_Dd%�
����S�m���o�×�+5��X}56�P�6��x��l�S�g���ɇ�� " O�����x܇�Qmb������?	��GF��C��p��K��כ�(1���<x%"/Ux&Gzl�+�.Uq߁�G"��;C���"�|���}:��V��
����|�@�5}�|����<���ͬI��rR����9���,3�?1���~�m�U5��eF���SH��bEh�1���2�7�VI+����9����U5�Ŀ�!������`����N`'��>�ȕQn���}�ܒÞ�<!���4��*wT|�����i�3p�'�)���O--�:�~��,m#Ft���T������, m;��L�8+jJ����J~���p��i���P
/
��T��0��QLȱ������x��g���/���M�&���[L6$27�t��$d�!��Pk��#�Zy��Bgm����U����M[�fee1ϖ�VK����b���WL�鰸*�)��cQĄ��Ųv�ѵ.�dD��´Z7�(d1�P������|.=˴Zp��G�:����z��6��������(*k�Mĺ��r��W�U�8����b�n�l �t��9T�x�X(�}pӔ���h`~��/6e a��	8tQf���>�_v�_zQ\ڳO�V`�@	v�ZE��.�r߀z��Y�DC�f���<��>���1Q�n*J	���P7�d�Í�B�%n����A����6�`�p*E���~���֡��0�(p����D�ur\�����s�
����o|�f|�+|!�9�ug�������ck�HXE��6J�N�Y��n�X�$�L��b��~�� �\�����e�[	�CF��� Ms�s���Af�*�X�S6o��UB��>{�/����N�e��wi�;=�m.?.�8뼽����G|&ksҫa���j�F3����>A�������A)W���:ٞ"@�e6��ec�'WHC K�A�s~{�����;/��|6��Ǟ�R,�]۴��#ִ� �F�>n	�%��rp����WM8��L�*��4~�-��2��~}�i>���(釁7K�Nuٙ����E�(���ȸ{b����x��CK7+3��	��J�Xs���`�q��GTN^0Wre��mL�Ԟ�����J�Q���^��]. n���q2�C��M��8d�hJ����ޯ��Y!�߷2��Gݩ�̌@�����=b��w(��}ʤ�-�&44�-�N$Oh��)�w�����|Q9n�k���nޓ/�#�)G�����.�脙��VCH�#-(�-��	�c�+�⮜����oznN�6���zV���z�[Jn���	7��	5��S[JW�'�2��|-�o`IVV�ҷ����5I6-���NP$�wo�ٻe�n��_�[P��^ȵ�`�0j �Y�B�R����VЄ1��3��ZX���	7%�
N϶HdQG/�m�����&%�wO��tRC�k1���A@��Q����N�h������y{���?�R̚%t��0�>����A�h�@f3֋w�G�B"��
��x��� �G�x����u@;��3t�P. ����T��� {�z�i����~��b�m��ۀ��B�n�U�_3���@bq�u�L$i��8 d�[�O��sq^�jMփ�s����oWnN�2�ɏW�Z���A��"��
Vu�ضeSkD��!�_�A)8g��s�+�hK�*g;Kۼ���#Sw�z;O�B�tT:4��?g�S&����H Z/2��v'o�g���C]$��un$���zܦ����,v]�d#s���V8�PN���u��s�B����������W�
�3/�������y�0&� �՚ˠ)	�kW��eB�΢�Ox�.��ФP���Zƴau�-u��D����D�r�Մ�ʔ�� :�~�)��`h�5*�d�E�I�b���(�u������vsRل��p{	9I��@u�;�Xw*�"g�^���xYD� b�q�t���~�]^x[�2�m����*\��l��+�Q筕AN�E�;�m�6�+.�9 �/�?x:ņ�4E�[Άȁ���W�(NG��/���A�>�1d����.�g�������d���F���+�n�2�y74l��������K�z�俋.��)8j訸���U�d�_�%	聯3�Ë\b�`ǚ�i�r����a�,jd�s�G^���6o4�΁�E��	�m#��x���d�.!	Ϛ�p��2�}�/��}�RhzJ����U�Y�|�͊+S�W���}G7���.3Ā�:K�o.6#)�x�=5�1�W&����ӂ��eF_�>Z)p�He ���»��Ѝ�HC���a��Mѣ�������}�w�,�� ��,��c?l7E{�-X��=DM�n�	C�;����<E�;����С{�l5
��5�	~t'�
z�b�oܷ�����o_
�V�mOC��@Y��y��F�0��)i���~��%����,0P�X׮����?�mw�&��߳����k{�z��^�(ޭ=����yG�7��)N9G���%���!8?RxW\�1���ya�M}{�����9eK��i>�eiO[��9�_3��@WOf�� �N5��E��è�iN�7t�Z$:?k��2��&�W��D8?�KF;���+�DH�_<�['���|>����L�N���B^�#��T~~ ��fHy<�DHL�&�M�R8D���,��T<H<�/����Si�͇���,�Üm��L��=�Qw��p|1\;�����6{���KEC���ِ�Qe?�o�Fkoo�X
B������i?b�C'�)��Q+j�u����ԁw7�+T&�S�7F&��ٿF������	4f��E�kS&�j$��A�د���n�u��u$&��Fk����=�d z�sbd��G�W[fd)[�IP�>�:�O�ůw�[�P�$#��r��_"�ax��&b���N�i6d�1^+%�Y�'/S�Bs�ߑU�_���)m�T\}�'&�x���]&4|�l��d&P����Ҍ"\J#N��6iN�
s�c(�o�(6}����gw��tրM�L�6�Ov�2�����H�/�s֡a���Æ��v�N��wC~�jC��������An@A脷�Ic�h���re��|RZh@�s%8j%�`�^���D+K�w�0'Aw@{�lBl����Oa�o�"��2ކ�?�aOqk��~�}��Z�!��Gg֙<�	\���D�)y�ѩ"�M�$�is�#T)]1K���2�cvW�p\i�]/~B�:2�1�����H��$�v�dM���q{mt�׌�ǘ�Bf��6�" ]�����)���hYm׿�a��Ԝ�q+vL�Ye�M�488�+ύ�1[n8I�Q�+�	<[�(o��߱f��gerC�":��.E�b\���ɞ,!�9 %n��o��~ji�j��Z��MC=���qYB�<z�w�ۘl'y�J�:��l�lOh�f���<�@2��Au�-��,����R[���Ae�t�"d�rx��'�����P�H��m+Ȓ��B��CQ^_e����^g!��G�BгD亾�	&�Op �	5=O��=�"1hu|׉A��f�c�]�H�u��Y�ɧ~%��۫i<]o��-�q}�5M,��5����¢r�{"��O�У�d7���/���_�viej�F�}��bq���2�R��r�'Vy�f�S�����(����vq������Q,n��)�{�C�5I���
���y�B��)��vV8{�#�_Į�SҊH���8븱ᰭUK���
�,aכ�`�v�.�R��+~�uX�?5`�VP���̑��!Pc)?�	�Hh�5���(���7��2A;�^o�
A�b����*�){j�'w��Q�${���&��E�����'A ��=����(����D��$����D#�o��%���9�}�*_�{���J\5%E�BH��$����[������g����>\:�;r<EV�R�Z�2[u］��O�k�q&�Ƿx�&*��,���sӾ�3�R��Ѿ�udh�KO ��!|3�5Ҭ��}�࿡��UE�|�
�J�kĈj���f-L����u�����8����m�6�6
B����<��I�VV�xӢ	���#�rs�/k#�f�k�R�{6��B6��W���u[�{k��ȯ㴵�2�����l���j7�3[,*�����%�!N����<�-�%ש�S�]S�$.�'��MMQ��Y�|X�.@Q���4ܖٔ��ũ�*6p��1��E��Os��#3U����<`{'�(��'�4`]�&���� V8CeXȷ0U����\&8|�]���W��ԡВ���6�M��E�Yv���ċt-�`s��L"@�!��"ڢn���I��tB(`')���l����Q=]0h?�����9���6��k����кv�Ї}�i��%��`���6�Y���k���%��/�k����J�����т[����r̆���1�3������Ӈ����f�%��kX�.��El��\;�,`�0ρ�q�iR�uEd�m(�B�����O��}}�"��-냘�+J�?6���9-t������cv���O[�u�f��I92(���(Ӳ��k�k}`{�WI��hmvE���!�O�p���r��$lB����I؄�^ �� ���-�Zm�ǡ?cW�ȹ�$ؕ��O����qt@��wcǞ@�i�]�P��M�5i����Ho�ӅY7�� ��[G�&3�<�ew泤�)L�{ ���οq�u�lS�>����pv��VR����d�)�4_O��RA���	a4vtu��51֜I��F������xg��5��㗓;̣<�3��kJ�G&K3�G��Yx3�IQE�.��7���5��'���%UX{��r~��v_�dڦNdYen�c��ձ�j^U��GK���)�}H���3�  ��U,'�H���E���$�G#��i�<��>�M~  �ra��w�ϰc���aD��Ƥ"�5O�ye����E�/;%5�'�ޗ}�
m+V$6>�,_�ey�6�Y�s�eNE�+��"�`��
N�?5.��j��3�PV_lKd*��r�Ơ;$?�6��Q�d�r'�g���y��O2d�B��"��,a��n�P,<�j�i�!�����ehX52���m-�f���3G=�!�Rk�3��d?	f�Ղt#��r�
}IMv0k[pM�r%h�����%a�r<ď&�qù��Q1�h# w�]�� v�Ge&֠*}��l���^���S��Z�������B[�����P�}�giI��]E�Ŕ\����_�S�hTst=g����Y�P��8���5�(�6��dؔנ��>�'����5C�C�O'g�Y~�zK�O�@k��]�x}So���m�{]k�B&�]����$�:�����~a�7�TB r,����{xIl�h�؀ǌ�ϼ���D:��HI�|�����9+7M�bM��-"l��.��}�=�2�%���7� 9=�]m}�a��Vׇ�\�f�:2x���"��Q{E���=���"}�$q��3��ЉQQU��u��k��c��T!�5~��N��/�P5=\i�Q}l?���*�h�]�� Aj�v��W�=�f��K��<1D_���֟>��$I����[c��T�|�JD\�?΂��ʩ�Z�E��"`���I�轲�T�f�&�L%1��;��Lt(]i2P�I��g,$OQ{�4��M�)>�\�O���߇���32�����%�@��ԟ����Jܳ��f;-p ���Q���s��v�C��30��<�ù�$�D4��K#�����xh�ą�6�
mW3�������~�V9כϔ?�����@�n��!�')E_�q=@]�Ġ~�)�2�����żE�׋�r��Ɣ8��2N◘��=.�D�	�"k8G��n�_�\�j "�J����'^gS��"��y�IY�nli���:E�}�2ƙ��\<�F��n�c��.�-��+��1Y�Ց!�p��fպ��X��:���	zg[�Cz͓���6$2ث��i��Չd����q���hOa����e��f�x�Yf�xYo/Ξ��O�Q�ؓ`��,^!1���1Qt}���:g�mH�*��Hlk��|����Ɣaj�]�g�ȖAN�W�M��\Y�0z~꺒��m�� ��� 4W�d=�=)`V.�����Ȓī���d�I��1��������o��Q��>n��Tj��/�z5�#(8��
�p���(���ه�"��
��e.��5���ǋ�Wi���;gR�}m���5y����+�;F��Q��w�$��,pC��ηvl�����Un���4���i�&�ATN��t�H-��N�9��o ]�͹y�g7a�JL����!�yh�_�ݍ���>���V����_A�$�B톫H�m�3n��;CD��	a)5Re9�����Q]���[dj��qP��s���86�L��D0�N˂w��b�E��d)���i��I���r���A~�	������- ��M�m�Q|^�o㭃��~�<�3M��8��=��:k|��r���4�Ŧ%W�I�~颶�Q#m�}�����Pb�*ߵ:�+R⥂�����h^9�����tw�E���S��q;3��:���������^�z�yB<Uա���+�D�dZ5��gEX~�8��iB��L7�L�J;����	��C��2���D	}�??i�D� ��ŏ�V��Y����ќE*�H�:�5�F�D�x�X7F����F�n�1(�������dw�@��8���r�.�"Ur���]�H7�s�#�r �V�9	�rt�$��$��QR��';��E�^Zk+Ļ��dC���˿W�9)a��^TKz���k��ImxG�i�-���7�>H;�sϱ�W�&��K�&��$��B����݀��+�>���$���`g{������1�o���mI�{��-�����l �Q�=�)/fg%�)	�+]���P{e(-WW�8
��jC�|�`Ar�����.���Gz�x���-nQV�~�^{:�V�j��5U�upMg��j�h�g�Q�W"�SJ�H�P��iz�sĹ�:��$�����e����p���I��"�m��&�,��;Op7`M����Y'�B�p��$��[���vD��O_�w�(�=��z�<?�E!y�]�.�B2�W9*e#��㉁5����<�U#H287\UD�Ǹuf��һ"�o<J��m��tJpU�	a�Y!<ao~t��Z�M��p�)E�އJt�H�?�ؙ��t ��n���ħs� s���Ә?WqXC10i!��o�,����-Y���c��^�]/e?������<�D.��O��RZԒ���|T��f���@��. T��?y7i{ƻ7Щ���#��HU8�8}}�uD��7XčJ�O�h$��Хh��J98Bs �B�U�́)Q�bE����]8��d�m!��X�uBr8�8m��W8p��1��n��o�`��$������c�K��"W��s5�(�f���h�K?���0��[8A�k	��@6��r|֤u�� F4�6|��a^dY/,��f�hs�������C_�tg�aϱ=P�.�sO�.�֝�ajU�
yM;�	�s��]����y��Rs.t�Γ�s y��	�xt/Vٶ���i�{�D��!�k/~�U��4f�25�0Z�q���7h�����9ݜ��<a��)	�1�G8��K�R�Bt�Y{%c�M-?y��S���p�E2ط�8!���{Ύ���҄RGǧ��E
2o�)xZ�z�Ϊ=/Ԩ������,ovZ�C|���Zj�F�����T�,��(gH���)�&bŎ�2�,���ӴOx�/x>�+Q�o��u%��G�9��߹R�]R��u}S�!�+�#��;Q}ޔ�3�7ls�0/������y嚑J�/�>���}5�0�W�b���P�x���~(�S�)���MY8�5��-�8��+H��\���]5�{F��...�ret��Q&�w�����M�e(�i0'�����]42 �ds�K�P�x8���l�j�U��ve���+�X~�<�zCա��۪ ����07��֧c����{\uHN2�ň�������@V�O�����"��ʳ%^e��'��#9�"�;�|,�lb��Ӗ�9)�ON���駏�n��?z��������q�P�>Ko��gF�6��d��n����6�"�C�� �	<���s��m��m�LkA	�q����,�����%����U]D�!+�g6�?��{��h�0�T������r&&%E�c�C5A�#�$�> ]�&��MF��6"1�Z@H�St�i�[����H��$,0�J�S��� Mp��J�d��,	�f���Q��k�I�\^�#�`j��ʊu�� ��}�X,��{P��S�4�&�^�N FH(��ٯ`Rs���"c7io��Q���F�-�I��>@�$	�*� y,�s� ��*˖h;����t~�����X�s)c��)|�y���xi����.��y���M8t��N�;�9%AȻIA�7Sg�`D�����=L��qj����X��3驀2f��ǿm��kaY[@F�0�F�R�=����S ��@Qu��&s|��w��N��ն��m��S^�:y��;�<n�4s�&~��b�� ��s��u���V��bK����9�	��&�"�:I�{+i�F�$t��h�Ya�~��1aX�_��-�ygii����?�k��X����b�'�]P����>
