��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�05O	0ol�$c!�@ʾ]�7����a�
Ms�����ɈT%'�u&1�K���w�C!:}�*����K�t13D�ӳ��J�|�
�(�2��;̠IAz!))�5��y�vA#Ȏ�6~/�4���I��i4_d꟞k�逸�f�N�uކU�J�c��n�)��!)��k��z��r�+��>�q��·A
%uγ�/�׈�8�4�2��l��:�n&ջV1��m/TBw���{��,�$�u�w��8��k�Qs�x.�'>����Ӓ-7���a���ok��>33:xV��*�j�o�W�W�X���p>a11��};C$}R]������i.ŋs�=�b�%3���}U���|<Ğb���D[�x�޺������5Y�mIU�n��A��c����vxZ��&�c1�hp7
/۳P�^^�^�����'���L,��w��s��
\I����Ic?�Ro��8I��s|�=�(����) &/�����c�'ݑ:߽s�,�)���<5��f��^y���U�+���Մ��ϚoE}!)��	>ntX$/�Bn���tY��zZ�m���f��尤���}c	���}ƺ/k:\���U3P$Mo� �"�]�j�n��ϣl�����c�^����`�i?zA�R�bq�"���c����=�Fm�a��c�J�t����	J'�c�$�j���@*5�ʃW�[�Ku�&眵;�F ��mp�l"�o)���o@�͊�ڎB@�`�z�ﵾ���o�G|�8_�e����Qñ�����!-Z��19\�7��9Xd�k�W̽��qy@�b���U����^V�~��\ҥxhhs��j�gG�2nL�vݴά�dy7��G3h_!�nl�s�ab�?�<��lJ��EP#01��2��E֮���+��J3��+�����i�A����ـ��,�.����@9���B9�Q�f��c�h���zj/K�����A���WO���� (n�V�_���£���
�lq�:�Ȍ�}���?>�-�HFC F�3�����)��J�H�-g5�6���.�����ߔS��"���񯅵����������}��sCy�~gS�ڤ���B�e{�H��gd���?�h�˜cr:X���o��:��^f�c���55�U�0w������ƍ_�������-�l���poYM$)1�Jr��
