��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s�����חW�#C�d�z6+9�@�I���@1qm{���W!S��%{�kS��x�`���&f����}h��˿�
xW�E����_@��{1�����G��%c|�����ث+22z�x�u�^�=꩓�?�^6`1dx4�W��^�>-��z�#�3
-k�o,
y�6����_�N�AO��-���0����r�ͭh�҈���ѻ#�-�����E�Dڤ?�����������i���ѝ��}��ϒ�C����vu�W������RT��~�:T驦�Pf����E �ܯΓ���f7����'n�F�:I�%]�b+���8$�1� i�J��.Y�Q�����֡(����e]�&�u'īa-J׀�H��lk�[�+�C�2���� h[�R�����rSM@P�yd��yU Q"(f���ВQ���]jx���\!p^
�yd����1����ߖjdy}�|5`8ݩ��RY�)�����߽�0��G���g����q������&D�!�����O���A\%u�{�sD, ���2�$�{�eC��D��t��p�㝨s}�qQg^��@����)ޡW�	�Vv�e�4W��$�oQC��QWA}���\����B+���� W&C,�ke)��(������+�Q�9\�3�܉<2��_�K�8�v�S"ˤ;cg�^*4�T�˅فhI���*,� o�\�e+�WLF�d	��:^�J���Y*��K��äe��0Nb9�%@�f��������` t��66"�U�6p||�nCf9���}l�1����wgk\;�<�.J������0Z�l���Pc|Q�-˚�l[ٲ@�e�p����Z�ɮ[J�w�k�K��XQk��e8${���IX�e���Z@��Ljp���w�_�u�'HU%��)�?��@��(
�˗�m�}PR�b�P���l@p����_�W>���i�X�n�ΙO7�:����$��znA�#h�ėr�G����=����i����R�@}'V��!]M��+�D�!F������{�sZ���q�'�:��o�����kK'gUC�ub��Gd_hZ�棺ٝ�/l�� {��W����$�_R�@��V6P��Q\�|�"��g�=�w_G0V�zzD�����FL���i��@I�֖s����։�������-˖)�^�\��EH�{�k+��u��WKBo������m��p.��Vr�=<u:A��F:��a�zյ><g@�WE5����0��)
��r�gv�<6���j��FЉ�Z�`�DBդ���DW�^e�rj�A�S�Q����q-�5!V�"Xק�ˉs�o4F���ﱄ��*3e~�_�vV�8���w�$�y"�#u${M8�kjiFM��ۋW|М�X'���fgm��#��R1�a�ϝ��- �8i���\q�l�<��)��(W�� �"�ћ-a�nR�6#�	��&c�5�+�dǟ�@舭�WO*;�`�ð~�`��B�� ��C�	�nir��g�[� }�z��\ퟢg�hQ[g�?y%�q���%v{9��L���~��w���PPݤ�N��k�0��"�{�7U�Z�Ss"�ֽ#���4�G�,H 蟤�DT��Q!;F$�,��A�|�ͤ65�ҫo�+o�V�V�`����أ��2�d<Y#TQM���K�N�1�}3|�����{���]ˇb����OL8�vY��Es�,0]�(�2��Q�Tj�%UQ, j�+��T$�pșz�78�fp���S�!qc���w��n��׫55M/)ԙR�m� й4N��}�R�M�o�.�}$_�<38\��DǨ�4}�a���2���#��O�_z��m�Fs\��+^��m{j��+P�ɦb�-��qZ��ۗ�P0U��}+��3B��AR�qQV�j{��tm}P�{�t�-~�F��W0�J�q!(k��
�*8Ȉq�>�P�Dw-��`�~�wXA�*ۥcS��3B�o�/7v���ni����1�BF���=���JPM�h]�z1e���Q�N S����N[�OKZ�:��\��q��3�}�Ǐ��Qh�'�)����Y��eĴ5y���҄'�#b�W�ǒ�N۾�\��r?������Գ�P�d��O+��i��lE�C�kXR�D�jbM�|��Av"$�I�,�@�Th+#\Y$'�Ci��������p��fW�_�2�f
©d��.N�gg�W|�(vb�K��pw�U�8q#gx;?�5�$,V�ï��V&S��<�M$��;;Q�h�V�Ao�Ak7k<X�}[8,{p�mAmD_a@�T�oo/K��]�~����к;�
_�2�A�V���c7��'K=�#o���,37��7H��v��J��+!��yz[-/��G��ݧ'3"�4H�J��U: -+����å9��x&�1��cI��/A�#FG��l�O�x��l��e�������/M� ��_��ٿ�`����)�Z�5�8�b���K�2UƁ�сħT2!0���C����j~v`��:T��rTי�s�}k��ӳ	$�[Ҫ
RK�0��Ӆ�~�reǻT�{����8�� ��	�3ɵD���-).~��Yc5~NJ�Y��Z�h�TY�M�L�r���Jn�S��|��0�������:h��GʥhɓD^��h_F��uGM<�s��Pӗ��#О%�@�Qúc��E�Q�IE�Q.ՀAꖏU���ɻaѶr���������#8KP��z5��z���Γ,���bI��:�ք�h9<o=��/�A����cAӏX�u�ɿ�Yq3��Μ�J��Sw�?U
8�Bhh��ú�1o�O�7nHZ�A���%�?�*]o����h���[Y��s����v<��l '��t��0	׏2�E�w��A��:de�j�w�z�
�9F�Y�5D������CBL7��)G$���#GQ�.��VG�\k�C`�-�$uh^��/J�֚�+��Mr��Y����@���ə��4+#����z����q6Y�d�:���|���a�{`y3��m��oj�c��)��@$����?��ba2�I'�'�:�����#��K[���ј�*�iP���պ��t��XP!��$�����.���qSIUGU�ժ�pj�O����Q����!w�8��i�;ȖK8��j�f�����2�����)Ͳ�JR�^�� إDm���M��.�*�j��!��	��5-����T����"B﮹ˌ��.��CD�j ����g���!�����;���,�)�@�n��� ��Ü�n�h��-���8�@f����m�J��xQ��8"W�G�p�D�&�q�S�4�*���X-�?���TM���V?ҩ��׋cRQ�4R[=`��y~�s�fz�=���rZ���OV(�D������'��O9'/D�T���q�B��(�T���l�ԗjĹ Wq|c3oI��0E�窒�jj�J[m�ء�"�*�'�]�x�8������G�ǝ�Ό�+��C��y��u��H���Ipcϙ��8��������@����u���Q�`>�'�
U��V/!<i �2���h�O��aܔ���>�g�i���xG%�=/�\���@<e��OG����qsv&g���R!�����w���5Ͻn�v��i9Q%ZjI����j�=�b4��Eq{�,Y���<B����|�ґH_� �UM.�ǟ5:v@�:�mr�f�nUe����t*y{$�&�p��oa&����>X�!b�5�U4sX����fS������|��&О,8����C�Zq����u�Ҫ�c�û�UдQ�B?h=�����ˋ����m^��}*�Ӣ�؁�W�FL��:~pVks�o��1��7���q�|M3�oNo�?}"�4�Ԕ1�_Q�3��{�Z��-�� k���N�6��訕�!�`��"�T^i�^�v�����C@��_�N{X�o�����xI�CxoO?�����$O0M=HT��V�^��B@S���lH�1)��Q�P�W� q��׫0��a0�����4��얢��Z ���cՉ/Af���P�Q�]�h�װ�#�`��	�Y	�.%���H����e-[�����2�����"i޸ �m�T����4�8ޡ�)�Krrc��f�G1��C�}b�BA�ߴ0_Ʋ��`�x��?S3:q=��d�׊�U�E�ɰ���
W<E��Y����LwݫR� �[�5���[�꣗��ҟ�3`6���M�	�.?V�#���1��MҫU�O�����N�#��dڧ��-�xv"�
����?���f���b[���vQ�Tm
�Cȍ�9U�d��`�?��k�]-��6���,��,�>�:���,U�XQ��Z��x��0�A�I��y�+�H���=�S�XV'gi�;�X2*���S�л���gGQA_����kZ�$[.�'����:s)d�^��[���v��̩P"kp�Z��?�������>�ف�w�GX�b�kԯin[i��d�����ϸ����a���֡}I3�@�s1�Uk&TǮ�Uq�hAYS��P> N�3Z!P+����Bg)a[��bi"?�d~��&�����W�N\�OJ�f��6���?}�&������m}����={C�2��uF'z���H�(�'��d�~Q���9�ߕ?��d�0̬���6���CJG�+�� �OŢ���1�;��CfC���O�l�[�4��w�Ifl�R�q(�"���
oL#.bD�W�,me�-pk}�����{=����yT�oCs��'�@<�^~=dhwI����
n��
�l��@{�8e�INH����*V���*v��* d���������ű�dda����yw�CK�'�%:|,�B���w��]P�L8�a��|�O!F���l���q��>����F��Ъ��.�hH�_,�Bԑ�Z��q���n*�t���#���-�����ea���U|Vl���+�uK��0"Kd�	og[*���ϼ�]%���d n(������2>��^��0�jU'C��,�8��]@� f��_@L����Ǵ�~����үƸ`�,X�^ͬ���Mp�M�ә+��S��1:� � �>*�79{ޤ�V�C�	C����Q	���Rk�73/)3Y���S�{�ְ:��/�g/9��"�^=;�U�v�A)�G�ƃ�W��j��G�� ���kIymaG������+��Jq����?���j�Mb�����è�ꮼ%�o�ˬ	���f�p@�9��F�~�4m�l}�����u4��f�DZ�5����VP�aka&��Z��xw}�����b�%��GJlR!��������);8}g+�R��-�O��v%V�b(}hײ���t��s���bݗ+I]�©�ڼ�L�'��=h����N�Qo��mq���r������~C^��nz���׭�f+Hf�\��� ��^F,Sej�}��M����؅�ڈ3���4��b���Iޠr"e��3���Sy����<s��-�U���xZ��ڜ'= I�M���]����Ԉ�����.(�E���.[�:c=�5��3�'u PT��^蓡IT�z��w��r���O�O�NV3���8*� ����|��\��wtC���H�,��HGJ��:�;c�QU����Y���0��¼^J�4�뗟�dC�.���qќ����F�:o\2a����ϥ�ծ�Z_�P�\��o2']���E�pU�����Ǳ�9.L���E�8�T1�s$R���;�ϳ�QO�j�g���k����Ps2u��V�c��k��5(�S ��S��2ju�� |�[C�/I�IJ�k1􆋘d���}/Τ�ݳ�{�͠�V�������j@�$�¦�P%)p����>R �	٨�'�u�竲8N��O ��h�T�#�(bЪ��,�uT6���"%ʄ,�#����Ӭ pnB3�g:��ZM��#)���8L��ID&t��,�Iz���p@3�2�hcT�ݖg��e؄�0���Ҭq��*ǧf��։���qlD�B��~���B�|���`c�/3"��t��tHBC�%�⣦$\���3�P��2�]&D� Dn�Zwo�du�[Ļ�|�D0�g�i�Ò��O�ݮya��2c Χ���V��R)҃�s��Rl�Ǥ�H$b>��\���):�
/�U<B� ����O��nF9hش��{�ŀe���S!;b�0�6Ƶ���5_7��l�u�f��U�=������߭Aɂ�/�O�	s�2Æ��&gV(��=CX&�_�JIe��{�ꉇ�ȔRB!��NS�%�E�a`"�.��ôX'��;��[?�E�*����,��Eįi��Wn/VE���Վ�36�a���t'��XΓj#�����>��Ζ��?A�X[��D�;�9!Q�zJI�t�F���h�:i&�e�/�-8���YS�j�4Yߞy2(P���b�O��4�e<(��6Z�zB��(c���X�����{ܓ2,�	���Pr��\�9�cq-�����m����#�	ן�Kf
vV���FܶWG܈���yJ<��)���/hIII��_��o&�'1�?p2�\�mրt��e-j?G,���|1��q�д���
�Y�THU�p�� �dӜg���
�hK�)��?ݥ+�o������8��dO{ʏ��G��6����6�:�l�8����4�49x!�'B81X���ډ-��[Q!�S#�������>�Q�r�n�:�r��}��������t�H@N���"��]�������O=�(��i���?=�*\&���m����TU٧�A�3����mD�W��`�(9"E�H��S�2\���8��^~�%�O���Zuѻ��"���E���^I�^�-�Ƿ�� �	z/ev9��o��9`XO�7D"P������P��w����}=�� ��E���X��M)�]J����YL5̀��K*����x��U��J�"���I�{�{A�Z�C��E]E�[��thG��12�p��������_��T	Ϛr#1y�T�?f��P`u�"��M��T����f)����L��-�BvQ�@��'�˿�+رM-�N  �`��Z�]p�kW���ϗ��nXb{�d���d.��&u�+��1[�9�$�e����?g�l��H4�-F�6R�>�����:��w�C����(�����
>����G��_�p�,svc��5n݇�5���OqpT��ٓ>L4Qi1m~Q�>X\��ctro�oa���E��P{��
��?��<���9�"�RE�P&�ꆺyT[�s�x��]T�n,8�$�2
3������4�����ƃ��eןU��/h�VZm��і����мr(���w���":���@��J�*�)W=�;�����Y�Aށ]�A?��fo�8����r2.O�+v�u򉢪�xfQ^�D�H��>�	\��$M�5��V�Ł�z���X��×p��n;�Nㄅ\��V�99�<�c&�]Ŧ����r�\η$30
��f�3�u[*� (D�U!�Js'�B��S���+��L�f���#�߫��<��Sـ���Z���CűT�c�?��9IS�8�R�EAr�_�oڈ$r�����ϧ��9����P~�-���tYjÛ7���t��
�����W�O\�u�c�� �iC.�0��z]�m��J���hs�!�I����D
o-�&i�SwP�����:�ԺtjC�C[�"F��ʁ��?|��%Uz�,���8�T���=ղ��DyB�ڜƘ�m�K�l���x�	 S�I_�Wz��)-4ܨ�9L����'OW�wG�1l���z�-V=Z�j��K����s!�	MX�";�kr����s#�o��=z���a�\%����@�]�2�ss���&������w�Ժ=��煢��+1��?�3�ϑ��Qp
��.�B5o�!wpV�+䴰�K�l-�՘�*��q�#�H~���uB<7��p9"%��)�s?s��~d���(\�.�&&��]�(�Xݥ�'g�4��,���������|��%����c���ɖ��;ʫ��T��4��_�+D��o�~�y�NLZO�v�'�1�i��hZ�|�LQ���S��>���v�x'���ьy�q|7�����h�7��7qWI[��q�&��h�S�Lx�Y�3h�F��4�6��g{�9
rz�ӣ��|:�'í~��<!o���:��hwY����O4���7�޸��œ���m�)�����)mkTF���M�oҿ��n~(e
>)��0{ٙ �.���"��<חR��g�*�"���q����h�;���#ش
fs���9�� �壢���J.��q��6��0J��՝�Tp�1c_Q��l����b ����F���A������OA�ڡ�z��u�a�0���X�6��>wK-��#�+v0F7��W�ԓ�Ax[���P,�dA)��N�I]-`�g�pd��H��څ�������ANO��4�'Hj(����b��_�-@Ǻ�6U�4��C-����	Z�\
{����Bl�'&ܩ=�.�{;F�^�k�Z�]҇�@��>Y��$z�����0_�-��\�f��eJJi"�ۺ�@��!��d ����u�]�����{���S�uO����C�,4CFIy>Z��:o��S1�jn=�h�JraG�&��$������gE�
��3�#�n�f����)q	���d�F�e)�K՟����C^��ǻ�B@��Q�=����_�.ۻ�M�N�n�d ?_������[Z_�\��F:��eVϷ����[��9�[_��;��gA�#f�>�o+����jP���v1����Ҝ����� %94絭20�+7w�ҁ��.���BQ �P���F�3�K;]=�X���/�yUNjc3f*�%��-�Z��,�B�3��vKiDqbi���V��~���+b ՠ2�C��d8��_�A)���7��\ǣ%�q�4���o�$����̫��l^ ��Z���Ө�w��o��u�4�M`Ĥ��b�j��ήs�0~���L���e��v�ޥʣaCƦ��Ν�l��+X��M���b�E��<J��Lq�x��)�'�Od�B,����n�ն��%�@��oIR#w�x`�^�b���$=�����}�<6��-P��l�4�DXI�xꏼh��r"�f˨�{;	����3����� #�Χ���b=G�5u��<99�W�G�lV,.��cG��k͚��(`~��e��f�NF�6���˴��,�&����D醳��_�a��q�Ύ<����M�$7!uS_�A>0������"@g�zE�Y�������/�_��_�0i*
��K���A0!��:5h<x��)�>[����^�(D��O̢���ף�����������n�� G#�z0�7N�<	�tR?���h�P/�zb�fC�N5ZR鏂0S1Z��$��u���<���}���'��c��!�cjIbta�
��E�*��,��.M$�$��� �����9�"��d憴{tm��8{�ܩnjZ��R�z��E���=Z0����$�tĔ@�����t��9y�����vq�?D}���,�q�*�f6MuSae�F�����{|�;�y��c� ܄:tS��$����dnp��F�Ӣ��y�A������!�2V�C���.�~ϲ��k�޿���uFc�c�|?�FS�)n,���� �iK������K@3mT�r�:^m�
�_$B��;�B?��\u�ZC�M�-���;�>ӣ(��@M!�ߛ�@fU
7����҉�$�0H6��^iW��'ibom���S���*�6rD�����J�X	A%<��?g�*柌��P��!���\��!#O���Bo���$���j��N�ù�dO[��9m��-�Y�_~����3����K�5�{�|��������O?�eM��9��4؏ta��Ou�L_�E֩ҏ�G��F���&�s&N�i��i���S^��xn0��I��j����:���Hu�i�qK�����82?;Iʓ�.�x4�iq3K`�[�
!8��O`��Mz̚�ܴ���":���7��f�I�Wç��.//��$�(w�HA�Ƶ#�o��6������L!�"'�̸jvN��i�/4�s�\T�#�!�/q�Pb��&M���%]��,o��'(�0��峖_�ټ�Ǡ�q�U�>Sv흶~��(���}�z�%�@}ÊH.��p������u�Ojl� � ��ǻ�Ķ����"'){�$�T<�}��UsQ�GC�\���C�.�G��El��z�ł�C*��w�[5�"\x���/b}�V`�����1���N9��CS�ô{˹����ߊ��`#�̧��|<(��������h�N�H�c���@�F�z6�#AƼ��ŧd�"��ʰ�h��K'ߊp�p�~%���Q��Dy�H �5όq�C��Z�l%4#�uE
Հ, �7$)�Ϋ3&�۳�q�����S#hj�H�IH���K�͇�AaRDyɑѽ�E(�H6�J�ע��I�tLK$���8	��j0�>\��T�螻N$)�UK/��j~7�0��B��[�4�'�WQ�)�"t��'9��;�}�tx�D_F��H��ғl�r��S]mnhnW]G߭��I[�΋���P򬜄瀁�灅�-:�� ��r��`�q^ ����\Xw�*o�ȩ<���/!�J�e�ʉ�_�N�1��������11���q}[)��`i/uD`�4����"vg'OS���k�D�mWckpz�.`���M�F��Z���t��F�,��Ei�w/���� �N�z���=X�u��@�\m�j�O+�����SC��2��v�X�N�A����)>ֱ|�/�$�s�f�H�>�wu�ۯ��~��@Jέ�Ü���:V��N3�3��I�ӌa���FCY��u)�nV:9v����-��Y�~�ʳ�(�U�+[����O*���vщ�KC�	..��	��X�l����h�0%�!P�<�WK����y�"�6`����8e�0 �<p��+��*6e����<)>��c���C1t�Y�o�����k�ce��������	��p� ��d;����}�[m'`���d������ktA��Ik^�ei�QuI�3��%���]�(���S�$>mU��2"�S���V.j�&����]ÚKWs���%<��4�RR�n�TZ���疩�erĭ)���a���2yrg����N���1+�e[�Hs���a~ky[�!\���o�:��RS���=�n�E��&K��uOզ.?#���#���#��D(Kk������6�3�%#��f�Dۅ,ܠ;H�o����\� �e;���֜5<a���$�p�<
�[9E���H��f�'�K ���L�Q��Rf��#cWY�+��R��q�']�]�'L��1kE��N�s*kE�q�f����`��$̧�"�?��!��?�P���z�b��N�f�����.�=>����&��(�̇0)�Jh?|`am<���d<�,ʬ�j�>j?:Q�3�eo�5�`�Pq��c�W�s��2=5��`�h��4�g����D����.u\Ŗ�'��G��z��غ
?i.���^ VF)�a�L^^T=:��O%F��4���E�u�W�DE�����V����x�b���tX��̒� �Y�`�wF�Pi O��(�����>y1�4L�=C�+�L�8׍�L�Ⱥ�f��H؆�8<��B�un���:�#*%���+��
���I���ፎj#<9;[C�[$��S�kƝ;9uV��������F��4��n ��F6��i�J��%�X���>��=��b}�႞>n�^�ޠ��R3 AQ��	(�L�c(
F��+�pc�N@ \������r淑b7����D/��-	��A���d�=дބ_��y�(b��}�uQ��X�h�?�]�Yk#�vY.ݜt
�<n�	�ߎe0t�%Ý�	�p�B�R�w�fp�0iǔ�r0H`&���b��4B��WҐ�5g)B���d�K�����J���G�"b~�J���Ds��fH�A0�>%��0�$eA��,���,�H�⊮�''6;��$���n�eNR�MU�l�Y"6�y�8��`�f����X�9H�#�$���f�I� ��B�bz��%�}ɿ�z�$�S�կ��ydi�I�bF�b�o������e�5�Yk����w78�)�E��_N�C���$��'����%v'ԖL,���.P#���q/
��RͿ��b��wF�ٛ�/��G�vFr�d7�'�����M�,32.]�%��R� ɷeX����<U͗��w�C�(U���2�U]�w�(K�,.!VN>��W��͸�pt�TԶ��L��L#�W��+��_�E	DJ��P�e��9�|e��DW,�Y�[�(Y"՟P��x�H9�hE�z�u(�}u��B�!R�g)�s� ��|,�6f� ���5� �u��N� ����V�~�aYk�#_˫�{lkL�3_��y9-�P�0�3��B�e	��6�Zt���h�\�a�_j�;�o=��c�{�S+Huf5�"�͍EJrWц�P�r΢�=��~P��k0[���wa������G]�����՜-�������$�ۺ��I���%G�D�qV�~�TO��E9���a��x��]d��
=0y�vQeUI�����~��K�=����#��p� Á��&�N�wCZ�2�����?`�a�ZV�b6���NFXO��ѷ-�@&Q$�Y/��ˊ�."h�> �T��B�3�b$�
�!>^j*�e�<�3�:gG�?0��o�#ϻ��P��IU�y�ղ`�z�)?P,�0��UG�t��AVaƽ�B����52�k�ZFK����5��a!1�K��|WE$'�9�1}m"�����&\!���'�J,�'�Y�Y���P��Ї�����w7�	s�6�|P !\���4��N�i@��]�4ڛ�T���,�r���B����u�Հ�V7"���_��x<�
Q5�^�(�R��kT����0F8���w)�&x�j'Mj��]�Is~�d{r�6n[<i>����(<���7B�mALځ�$'����D��I-G(�!9��W�;� M��� ���E,�LG�&��k�S��q�Z6��te�����`7�P�=�l�aQ)�D�cW�*>���A%��,�!&@� = �W��ɣ�,��5�<�����c�E�j�]^䭨�Q6 �d� �<�A�[1�&F���'iY�/���oI}��J�{���-��d�m4E�r�[f�w�X7bU��0Gw��}~ɨ�}h`���N�~�h�[��h`	w&}��>�N�jD��.1�XH��O�����ÔQ��1b�p2�ᨀ�*u���l�(#3�s�Y]�\����w~�����6b�Bd���?q�{�%��?��ի�hO	+�Ȱ�F�����u+t%�f��	�U��Ϊo��dT:���,��d�Si:�O�Ƨ�U�8�>�f�rIJ�����$�'*��lHg�t�Y^#9�ֱ��Փ�����"T�?RON���9ڂ"�T�j�ʿ��/=���<���kHyqeM��gW?Q�dΦVӇ����k�C9� ��oI}���)� ��Tכ3�Pz��U6	���>�2��ٞ�/�#��E�L��1v�s`_u�V�H��FƹӻK1�/�R<���k/<����`8C�%CH%�����Q^��VQ����]v���xĥ|�T��P�z�4]���P������:�~���I�yw������P�5h��A��k
�]���3�ߍ&�&� �I��S��A�K��	}}B���Z�p5����6�$��v�wl� J��N�~1��g�g}!Z#�!�|�A:��2�=�p��r�P�1�U@�};X%«
��:6 �]���+��_�ُmnZ"h6��ӗ q�i�K�=p�@�^%k�ٯ�� <:V�pN4[�r�Z�B ��h�gsC���W�b2e�����F0�]���|Fa��^'׮Nbk[˛cFᆂ����F1�'�齀�����(�7K���h�NK�dmr�I�=��${oS!x���T BXC��,`�.��WB���zsվ�odؗn�qKoJ��o_��_����Ӌ>t����5��
�)i^�$��k���4k�M]��mLg'���y�1_�=6w�i2fyS��4Nr�WJ3M��N5��<�G��g�}�oyUB�^�u�m��V��{����je��.گJ=�ܖ�%��M����r�H]�E\!B�	+�L���8�yMS�f�X�ٙ	�I	D^��!%� ��.)����#�{+#U��u�J�*!Oe�_�W� k5x4i�&>���K&���E�6>�yL�.��	�F`NM�%P7P��w�}�k��5�hUPr���h�]��"	���n`��V>Iڷc�^g����c���}���&U�qk�=��;_Ȱ�9�QؚR�O�9�Uh9&.�e�ĸlz�T�[��*��{́�����_���٫�D��(Qu����x�(.��V�.��6U �<�l��A ���K��k=����V��>����>�SN��G�h��e=�0�I���YG�^��!h+��BA�1τ���7!p3h1�l�z�0p��2�P�����(6���^Bv׉���l�����{�#Y&�J�LP"Ğ�Smv�'d���}�Ѽ?��mC&+5Y
)1
�u��Tw�v�"w��@CJ��������qW[,k޴F����!�E�f �DA��e���މ.�3�1Z~�$L��k�\���-$=��\��e�dﬂ��O\�R�ᒼ��W��7�������Dg���(H9���0�hЭɦ�?blH�;GF��sdF$�q�0F�fB���ۦ%�Qb���X���l7��
LXn*�7y*�֎3�5��1��zvM�o�qXm��ě�f]3N���㷏:�{�mC,m*r��;��H�� ;WF��ڶ�����Q����f�����)�|��0 �����k�r�+Sa-]o�x�`,��|��.;�����>,jϋNr r.�Zƛ]��.��C\��U������u�`�p�+>�$�`�p��C������9��`�N��q��}�G<�̓�@C\'�����j:��3rYc;T�_�%Cz�~�78��.�.�_T���c����1���x~+X@5�o��׍����(�<��k�Jp<[�`��5I��d�v�ƫ^��<s�����*�[��鱣����>*�c�(`(�73�8�$���3��6s�	@/i����s��$F?ѰDŲ2�WB��0&��r[����/�B���܃Ơ/1���aƯ��'�6ta�E�j��.|s�q��h㬺��x�s3`��~�'��	tf��͵)��H��e�@.A��0�+WZ�	&��˳U�%i�[�ȅ∦�Luë�I�g�0.h�oo�4����2��`Q�g���j)�h�>F��H�#��d1�党@�*^���A��\���!$���Orn�G��fd�[|���-7�ԪeV�v�Ah1���m�7d(�dV�#���C�/)�3Vu��f����w!Ɋ�ir�t�9��QJ"�E��~��2�E䋌%�{:]�i�#_>�2�ed%�F�Aa'��ˏ^�5�h��Գ�)4e�0pG�G��/+�&,Udwt��%���4֢����(^�BO�C�I�0��J��Dp��o��n('/�|]����r��_��[Y����u���׈��qa�g3����ᇈ�Z��+�BZZ�iuG�^_? }A�5<������ّ�o(�Y�G�fq�HV�촛t
��AR81��P0��i�Ēׯ�K�6�k��Y�9��s�H����y_;eT�ѣ�o�����u����:B���W4����Pgτ���\P��i���&���P;�8�nV=����JM{ǡSs{��B!r�o����P�����EE�2�����E<[?s���n���������rj�{&gAr�P�3Ú �YW�^���DЖp�/���A=��O��r��*�����Ȃ"��:��[:�A+���q�/0����#!�"�,>7w�ϭ�]ʃ:��P��Y5����or�5�%^c����L#�qWE�iI�k��x��C=s5�M��]��ǨT���Y�D�̸Z +-�G>�L�r��N�4ѳ�#�9�� �Û	L�Kw6z����U-�n�N�yZV�r�m�N ����N�#yݷ�J?zF/ ���<��u�ED}	7��AK��M���;�|`y3���,{|�3Y��%���70�u7sJ��؟8lS��a�P��fl%�Y�%�Ó���B0EmV���g8�af�_͕����y�Y<�� ���Dû5Z<�R{�g���q��P��ڴ��T��E��
�D��	�Q]ti0XЫ����<����"]������Ҽ�H
Q��_�VI}%_sz,ݬ��Tw*�*�0� ���Nz傼x��n �/%����(O����4���Q�$�)�b(��6[K�-��X�-a I಺T"["_x*8E������a���R�H3�ފ�\K}Y�����(n)��\@� �Wo�&��,
Wh/+�c��}ڡ��@[-׽""t�GQe�&��.`H�c����^��[}�riAF�	�G[�Y���x:'@��S�#��s.7��O�L��\��yl���Jf'���+�å��;�QA�I���Q�-�����ݭ�ޮ=nT����!^�;]�^ǑFW�N�����jj�g�wOPp�m�B3Ft ��f���H�C\������8_ ��At����8�.��]{K�PcXq�U 9l�����*}�"�mzk����l��H���@\��=dMS�h�U�0���ch�| ���χeX$~h�Sl|��Xx9��F�C���Af���svQ���6ʃ��[n٘����F:�٪{)����}�'tL�82&��V�B�--���a�t&�G&�=U���4��W5�;��۟.�!y�GяԷ�c��|�g�C u��o���;d_ohLך}7���>�Zʆ��p��[R�c���n��[�w^%$�W��7t�e-E�v#�(^��zC.�8�����q���o��	�ݴ,�!����4� �H���d<7����m[Gb*�e�a�)��]�tHoG���\��ޙK%֟���t�s��X��.Q��ߒ�UX,i̒5�� �{��B���e�^��+�֒��V�����L�����j~��oP�Nr)2����f����{��%��.�?A�x�2�ۻӧ 9�O�Z˘X��\^IڨB������`�
YDoy��K״?�i�TS7���4v�������>C�O���4!�@T/���EǛ���.��O~L��.���|W���I'�����Pu� ��=�w���	%��5��kU�	)�������T�Y�
�o��ۍ!GPs?e���f�<sӐ�����S��*-_�4$�
ļ�.z�"��E�5��ԋ�D�)����6&����1 �"�)g��iC�$��~�5AA����</T0��*.�������v ���%�w;��w�l�u�]�����1a���(ȿ��D�w'�M���JcR�mI�[�=ڠ��)v�%՞Tن��l�R{�B�K)r�*�w-�����g���_�{K��;��9ڞe (���oSNS���CTL��"�F�U޹���fF o7#p�)�Ւ	A�%���Vܝ"y+d1��G��c��T�Ԓ�F��Bk(�+҅�{�D�a
�"I|<�dy6<�uP>_��Iu/H&t�X�Z���le� F������U��ܶ��(��]G�#<��5W*}�W��Ko�ٖ}[��l͞W��Nڍ���I��LJry''0>��%dF.��"��OWz�&�ߊ(C-on(��qj�з�bYs�=9ln��ȿ��ՒD�̪��	B���Z���2Y��y�����t0�f U������+ڳV�dF�SH�~��G�*#�]�U�.�
�*fF�Z������1~�h{�}ۭk�A9�<�P��_�vD��{�nF:WL�4Ws>�mй�5�M�p�o�sZ^X�F��=�o�[�-XJ�"&���3UI>�@/�a ���M[�W���<ŧ�s�E�����єE^�^�YKP�$���Qa2ʦ��u6i��������r�հmjfaiY�O�CW�Ke����?����3LR�j$�/����=(�1f7[%@؏7���އ3MG�"þ�y���1�@�w��9s�`�x82� e6�N+�V�~��еir��Q�;�����!K�Cy8&^��r�R� Nm���ld�H̸	�l���B1oB��f"n�p I)�H�=����s�-�!�gfAZ,�4ֻ�[a�|��w�I��:WV0�J �fؓ5FaT�˯4_9�������0X�L�Zw��F���T�
�ǎĕ�AX��	}<��V���&�
%K�5.��������|�/��^��E8)D_��!���j�!2�ju�[�FV�`�E,#�JkN1���X�/5�ݱrM���h�9K�Q�J���q��M�X����lAn�[$uW؞Kk�1 BA؊ �%dw�8q�l�+8v�@Na~��ɉ��q@%g>äg�b���<��)�y)�v0PT^}���K2.�$�{��%H�2 �����@�x&�ւ�E/�#�Y������၊#W8�Z�6/�gۧ�B���l�V�~��:H6��7��Es���5p�?�w���,��WC����|"�J}�OFT�&�~k-Q6;��^+u�����_�@��lL�??�[��L^�7N�.Z��vkA���=�7�W,~��BW����-A�ϊ�׃TI��U�������:�Y��YEm%��<�W[`�6��̸��]z#a�
t��^�A��&D>�Zɮ����kcZwp�Ǡ�Q�6�uM֟4p�j䪟=q�g�+�X�ʱ5@��������sH�ّ��qɦ��'��D����g��I�`Sy͘m���1�Y�
r�����&����c,���o�pJ6}��	s<+ 	��m�Z��m4hc5��֥4�#e�? "	�2p��j|���4���Z��:g�?�e�# �B�	��|	����C��&��l�:ȴe���7�5����6�G��Pz��-�Z���Җ7��%v��A��qBO���j=#�I"��t0�rޘi ��˶�������8fZ�y�J�7�Q�[����j���5��C| w+c <��g'�V�	ݍϑ*+��
�p �z>SCe�~�V��n�����ᡱi8+���%a�b�'�2�naАP�n���^����C�K��i�V݃x}(�啃ǑI�_I���C�vNJ�Y��R��?Ro#>�2f���>#�4�&�7gLL�S��ԟ���BnV�d�Q��$d1T��=�͌D��w$M��$:?_UM,pt�L-{:d뚢v�cr�ֳ"�e���k�i.�()�)e#���ż��:5������		�rK�"��`F����8"A�B �;��&'I��g�ӊ��e�Epu[{��GoI�����ߩ\�
���Rފ�P�#z�)1 �n�D��Wþ�W+��-����_��ۈ��ǖ��
_D�K$��q{;I'n�$���ڨ���V>��R�[��;��2���<���f4��XX}���/m!�v���X �vYb��C�v�Ji-���v�,<��(�A��4m(��9�X�N�b>���K��W�*$fڇK�}�<q0�EiQc��U���|�������T�E�j�q����Ԛ�+���m����%���ވ�H��.��\7�y�H��)_��p�ӱv�j6)�s��5�Q��4�[�&�sZF��k�ۨ��9+���WLr��i�>����d�`;�8�&���T�f��[��<���#t����"[GM���哸]2���J2�џr�Ҏ�����'%�Ç���`�Ԫ��l�-�6.7p���9ױ�j��P��H��F�3�����?X�`��P�ڰS���b
�5�!��P���^TS���9�!��HU��L-�r�%��&����ˣL���������˹U�zL�h8��i�����e�٭�43G�R�IOG�ޖ�k<W�ln`\��WՋc�H�M��[`��	��s~qlu���^���)bSn��5�-d:���_ض�'��]��x�}�����ېR���i�C�7)/JF��4�X=�Y�*�61�%~���x������M~���G���|}9�D����$0:ԭ�O���V~J�rd3?+�$����T�Id��4���B��n����y�#�v����|85(e�{�e�Gw�Ñ�Y������T,O��J�L�k��m��͉���曡��n��HUs�*�Q�lt	�דw�O^j�R���O��;p��Z�@)}<�pQ�˴7�e��zS��{J�Z�Ё���'�%Z�$%�D �:�xb����fOZ��0#Iތw�v6sb"狰�h���jƌG����C�h%����� �t=F1:f��A�'`�i��orCE��d#��`���Qk���ί����1��yX���̗V9v��%ә��<,�ut���b��i &�\�;v��#�3,��w���?{?�rFX���A�i��ŵR���l�5m�!|�]��>�ܑ�pZ�|�RJ���'�֢n��!a8��/��$��@��\�Kj<~5��Ĕ�	Q ����V�T37
�S�}.�.U��\�-�nY�0i�]G$9�7$����*^"&��`���-jq���t4}њ[R�oy���Jv�
>�R��lF̀}�<��)3X�=F"���H�����D���m=C�No���'��	�9D��`n�س6l�Lt$ �+��3b����h���8(����,O]�T��z\�@v���2I��PWB��$KJ���kM&;"gO��2K���K$������9,���J!aR����ppS���\B�,ʢ';ly�P�Hڒs��('P�gW�C/��УiM�L	��I�R�?˖�	��7���sGƲ�l�C�jB�x�����:,��n�d�>
Vw���6�-?��ނ��v�0=�eu�N4��G���V���D�(����;28����z��K�����ß�P�7C(��mF�F��:׍ECT�y��� ln��_d_ Ƈ6�$�����"�����K>
=��o:�	��f�i��8�ʹ� .~��-�P�Ϻ�,�lт����bC:y��U
q���Ctee��s��cҵv��H9�����'�L�&H2_�=B�%�	���%8����~�y�X����t�	0 B�~H87��`R*�t(��7�n���13W T��3�^�޺qn��VeQ^�0W,tvɬ7$�DB�h"ש˖x�9i�<9��e��c�� ���;W�����
�]0�N�%D�����D�1R�w�4r��f�������G�~����PwИ�"��2�Xp��g������~���9�����~�^��;ٟ본������}���W���~Q"����y� o�`Ê��2��}��P�2����	���f6D�wڀ����^�9���Cρ��A� ���ch�����*�I�1� ^7i	�PV�?�0($%'�g�C���_C�fS����L̳�כ:l���<�C�х�S�ɏ���	�E�b��5�K������׾�[l����T�k'�s7��v��cZ�E-UG��ʖ��IgNM�O8�^�����Z�7 v+|�[�R�
�~fa��:�VP��/���\Z���N���q/bU��8_��w��/�go�/��Z�� !N�r�F���D4I�]�s�t�.��2�ן�z����0u~ό��dg %��Vv��KK.���ƶ�G��_l(���R�A���'�4�E!�!�s���1��͔ӵ����^^	ef $�c�k�E|�@vJ��⃟U��mVw�w~�Z�;�4A����Q}����G�� �X��e�H�v�)��=��t���SG��c	�W2�Gv�2T/刀�=��m��1� 
���^�q�ȋC�\��X�B�^�4��P@6�R�y4i
ފ>��$U*�i(��3�b�P���
��U(6�J`��:�ShiB
�dn?�]Iϗ�r�4W$��[��[��~������/Rk>�1���c��O�>�Rl��b*��_�n�=1oB\S��h�t��u7���חl�ʉ<���J:�0x���$�V3��72�y�`��rN�p,����6g EE+�6P�P3	��vƹ�6+����̆>��;J=�������м�ұuZ�A7�t󺠗ɻh�	����J��%A�>B��2w�H�5B��(�!s����c:�c;"0�z��T��GF�Ə+�ڿP�}�&C^fZV2:��?����H�ȹ�]����ǌ�� ��0����݋�O�ۿd��&�lfՏ0�L��j��}��	��,���E����1C������$4cFw�iD�B����啨F>@_u`]�b$������Z��)�x�@O��膹����Q���R���^�@�������Qw���pd�xw����7iြ����;�}�k���ɰ��Aኧ��\�P8���c\$N ���<�⭸4!Ն�gT;����]���R�F?�Z�&ո��ͱ�j%��e��k�Q1����t\�U���R�X(�	Ȅ.�{�b���`
�݆���s͊ ��_�s��Y�_?��!s}�0�o ��A��3�{�!^ݱ�M�'�K[\&��Lp��+�	�cc���P3:����t���e������l�ي����D���7�-�f�".���-�Y�Y���������d6�\ֱ�v�~�#���	C���ku5T���i�BJ%���ǥ�D�W攷#��=D4ֳ\����`z^��kz����.d#�E4x�����!�����X�n�6X��߻
e��eB�Ρ�sD�����6������O�;�W����ɚtJ����c��G�_^�������Zl���xK!�Y�Ð� ����L)2Wc=���8�?~�ᎊ^&�_d�Ȳex�-�Ȓ�0�]i=���1Z���&T�QGI�]������ �Tv%ȟ�*m�xW��P@qև&$�����9�M ;BO1{I�}�Imݢd�qy���a�[|���v'QVL=o	Su�
x��󕹾��X�3����థ�[k��l����y�t~4n�/r�p���J���D(��Yr�k���ƿF�<�������	��,8\���C���벯�&0$8	Z��"����M���H	�Fo�����?,�^�i1]}��uw4��ܪ΍��ʬ�
���r��#l�����Cj<V�n4Xi<�����|�F�ư��F��䘰��y�UN*g���zh����F�݀b!�#݆ -�Q0O]�r��iXA�( �݇Kc�$��KG�e#���[O��]yJ����1��\�?�:�$��%�G������c��,����\s��h�9U] ���>)�7�v���Uಁ��P|X����m���MǱ(4�|"�,��DD���S'��Z�(:�e�t����X@0����s�s�
4�}v��@�a� 	p**��~�Y}�}͒ᆚ�8� }*���if�a��-�2J��(�1�B_�0؎=]��v�P� Փ�8�V>�/�٬OU[Q��!���XfE��|��@�s�H���УFO�"�<�f	��޼j�h��T���݈��>5�����V�5,/�����+n�
�镯=�aRZ|�{�(1J`m J0zO�����Q-H�y��:f�C�ǁ�0d�xI)e���4�70R�-fy���i^B2�������"��U�-����©2h{��ڒ-h��|�e�S�.0H67N&����dR��2D��Zb��9�����p3��6U�����~��t�W���2�ը�E������.8�n�lg�\e(�6���:��,��:>�n���E�M��l���r ��F��^Q���E'%�h:�OPk�Y�d�v���7� 6xH+���� T9�8������	@ړ���QC�"�H��YlkzKq!�ۢ[,�"�#Z�?������I^�CŎǱ���Ȝگ�ډ>��C��~����k��M�U~��2x�p_�-R�:*���ĸ�^	ck��T�R�dAU��C����e���B�0ڝ��Q� �3D��r,�p�MѪ�u�Tap)�!iКƸ�q����_s&?���>El��L}��swX=����x�)^��cB���W�1.@yľ4�	�Yjh	�R��S�l��a�E
�~
8,̰{Z�k��<��/��e��(���H�ƨ[j�z8���3,��wH�`أ�r���B
N�5��� ��=%*E�`�j��^����zr�|��f�!���xi�-�r�0�����C����h�����!��fyi��j�Iݙ`�~.&5E���#A(�{�I��c�0v���0��T�bV(劐�|"����b�*�w���DU^F����:6NU8�k}S��}|A�5�������~=	P�I-�Ab@����8��xjk7jx6wh��Y(IP��/0f0eĝ����@�0Ѱ���t.�U"u�Z�7/�Y#�I����j~h=��;�v��0��0�q�~����Vd-�1+�ȶ�V�$�|�mOT�d��]�iR��>V���m�4�4��'mS}*d%�4����h���=_uB,ҁ��*RkjuY�����db�t!H��Wce�-hL�{����~#�z�Q'�J��6g���H�狞 �&ϔ�c���?W� ����~H������[PA˅m��2ݳ��Y�Jx*:��'�>�+��87D��mcn�p�u��($BRL�/&���C3��y��C���獠,�U8���xĽ�ޥ%�O�y���_���*W�p�$�ͧ�`.8�~T����F��z�C�ÓR�jo�M`	��ֲH�xZ��J}!�� ��4�[����Db5�=b퀮�|r�>-q��Z����)�V����2�4z�cC��;��V�4���fa��.�:�c)��6l�ݯ@�%.m}�ۢ��=~����Rɽ$���[���T�0�pȃ���aQ��c ���T@�ͭ 5ڼD;{<�̬���;������)Z��7��KW��L0��r�I���X	��8����ĕ`˖�rܡ�!���oq̝NP$���a�l�=W,Ɏ��X=V���$�	*vH��ּ4$�������0�Kgo�okq�6��{�����u����3B0��h��d
�w��r�c�/��#F��C��#��4�E{T;��;M�CL-��*l/К�;^>RRI�n�;p����y(�n��T�
溄W�݈���to&� �
����쒣�-��6!��x�$��v4N�]����Ǜ��۔+r��c'�̉V���Q:���&bc���8EZ��o���� �˛r�&%%����,����Q4����Ǉ��*kxP�W=���m!#�u����/W���s�[�;������ >&�*w���&wIvpJ�r����$��	bY��0~���b��ei��^��^��1�B��=������I,�pއ�eT��;;�2{��G;��X�|�d�*sC��r�UQp��Cߨ��;��{�H����\�H: X"���ؗ�`�9��),���@#�	��AG�k�?|F�Oɑ�R���	MV�+Od�؄;���ܙ�HqM����f\���7��oeo��Z�M-[�6mC�xJ�͢#���8��0�W�H�Aw׀��8�;C��!��^�L��^�i�ٖ'��Jߺ�r@�v�R����ʫR��C�L�p�)4y�^$�U(Y�w�*J͹Z���[3�I�0���6�)��J#����-e3����Y���~�5�K�p&���;HX�RU#���ˎm,�Qb��>>#*�����vb�5�f^���9R�yUI����˞�B4�B�����k��SC"oLx�'�i��iP�ͭ(
�ǜ����[�I�YyͭE���٩����oɯ�TJ��/;tk�������x��ˉc�����[�^q˲��܇�Yq�Zȣ�y���˟M8��Uߗ���<�J
Al�wU�����~�y�A�<3��{���Њo$�=ۦ�>"5C(��uwU�(�Q!6ME�3p�*����=��R?4ZW'R�8
�.1r`)F����g@�����Q~:
�/��a7���o��
��q��*�5t�S�[�R��Ȅ�z	�nDS�6趧�����ｎ,ob������˫:���/���?���ʮsPWuƊb��@��g#��*$�0*K/ �R��+��8���NE
w����;O��Sp���¾]�Y7X�� Z�"���JBW���5�4-�~�>�ұ�'9��t�Z%v�|�j!􁱹dQd>�g�
sU1����DA��a�Tz=(��ȍ	��G�4�l _w6����P7��/v��Y���֒Ӊr�F�"Y�ee %Ws:���e��b�Ga��ڊ����;�]Hv�^�O#;5H*��jŪ��M��QE=� ~�L07����x�*9W���r�K���6&t��Ք�˖���~��p2�d��!���rx��*�o�h&ÖE/^N#&��gQ:/��d��ZIP�.�_I�Z(�Gs7�N�Ž�Z:Y��h^Zh�:��q��v������_b��1^�YpiW;�Ť����w]��A�-ĩ��Ƃ�4�:�?̓�R���Z&R�zn=��_���C�ӄG��hz�Ɍ������
�ِ��-ȩ!1ai/�r��r���W���2��f���b�G�b�Y^�jh<����d&1��n+��Pa3a�YL��%V�L�q�Š�ˋ#'�,Ǉ���7����+��u ��� ��(b���rF[m� �x;\�@����j[����²�l���j���!���D��v^�Vw#�\,Je��,�Y����FFY�ט��v�4�U��;A�:��p�w���|P�"��wj����. ���,e��[v$Y��Z3�
���W�����y�L�alg�_HR�9��X��+�O@��H1}�"�@3 �Q?��� O��p�_�x��B�?����(�����Mc�%IMz�����-��x?��#XR=z>��X��K������c�P�	���h��Fz0O�ްI��E��h24����\���G
6��J�a��8�z2)`���?d|��	�� ���c� ܫ�H�mWM�m�����51���������*����]3X�؊����B��0�=����=�hk G�Xa]C]��+�&�X �B�$������V���?7wF��cZ� �SA�3c�|<���񊈸��aGD�5m}���U���>A����ƅ@�N��X���r����� ��g&;�sk�f�+C����|�6���A=�@��F8��P�m�����03�ـf�)�'��p�(}��$��U��=�V�@%���M�����JI����8��|�^HT@Jp��WC�Ae�+G��0��s�����d���-���֔q�8�&�wB[tT�Z�w�L$f�,�>p�l��'��g���y;��op�-�Kb�nFd�&���*�z�����g��Z�G���IGƻ�Y����}�c-�]
m�	�,:� �P̒M�Z<���?E�5-t;	��
��r:�����|�'��<�W�Q�J?N>2X��{y�<L��o���Z�\RC��(,��иݠ'�%e8*M���p?��*��6S6���)g���{	�K������13H(ֆL�k���(}���zuݐ7Ji9Ղ��|"8n5Gjq���O�� ����;hFf�]? 35R�6�
���u'VhٛGA�U���e�bȍ����c�(�zFG�� �y���V� a���G]���0��!�����	�-�=W��G��	�D29ƥ6��['�˼����-�,N"ϊ�=�°���k%�Bc��Gdo<��G�⚒���;�f��蟪5�q+��T��o~�,s�>o�'���'+T^'[�4�V��|�<�f����`s�k #}��.i�OM%��ed;R�؀;d�sӓk`��c-���+we��a��F�5#���·5^�dD�F&���L���3.*u�AY��]n����Ņ��.��-�q����eJ�����Q��s#����s��*ȁ/N�R�ŉ��U�yh��$�S>�FL9л눡�D�U��Fy���.?I�e��PzY1��8��RP�/Ou~M�������U�ù9�:f+�$�Cο���=tZ@	?r��t8Ӓ�T����_�*����(M�JG�G��
X��{%u #02)�nx����U{ ���t�i`IϜ3F_����KHm���
�R\�B�M��J�T�u�g�do,��sO@����6�fn��=P�էoT�aBy�+�Q����'��]QG[4�5>Nf[�����CV 9RF��@`�ֿR�,yB��e��Xh�7i�n:�	�[���M��5^%'�(�~�����?$ue7τkI��5H�]�L���׽|���"G��{�i�
w����ԜO�">��s[�Q��랂K��UW�S}�I'ϥ~�Lz7�f��`5���-ɕ{]k��F^�[�J(��䁐'k.�Q���͔���:��-�$s�aԘ�H����L��M;JT�qk��s����p^�(����)ܪy+a3�"��h%���MwC�	d�)��U�����z�[W�b����SC;YZ<)�)m���o���|n��3G,�o!�7P�Ê�_��=��(�@&i��wz���/����O	Ρˌ=�z��)m�Z��Dbc���tg�]�����1�HntsYlc5��]��j^	���u~|㹸�i0�d6��c��0_^������qJ����r�k�<�҄��ͮ�EXg�{�n�M0� A���x�hp+�M?�GixԱg���ۆ��%ď�/6'�®J���*��y�^�^ڟ��awCPO��%�g� �ԄQM�G��01�)d��b�+z>ri�&�\/�h\�>��J�F~F|�?Gz�6OĿ��r��6QL5u@�/*^�SZ�vԬ�x��:�<�[@?3aln��Kdx�B ��/�J}� 4Z�3A��
7m^�M�s��:Vp}Q���,�P<�]�u�F��_��ن��`L7�7zd��@v�#-�"M*G�O�ؒ�*��ĤI{��/�
"{DY{��Rne��	z��zE�(Hzd�V�t@f��\w,u���vD`pӐ�{�5�ԧ���a��@.�) uNH*$d�E�`�_ߦ������
m͕.��:bl�0��5����3s�hAx�f���Q'a���H9k7�P)eqʇͽ,j��J|���zL�����uoV�0�ǀ��.h�aX#���/9��F�v��j�)�����S�%�������s�T�Z�w	�[܂G<F��0�Th
/c搝�@�%YF�i�Tl�Q����U��8��Pj��̍Ylh�e�����I}p����k�8�3N��羶5RiW&AZͻ�M�@ǂ��o���[O�gB�����u��`*?N�h��`�������ZG����T���q�\��a����m�8B�I�C,k�fE� A�{��Wic�Ӝ[�l`��s(eڒ3�mD첑3h+�x:�f1n}�jm#|�,ƉB*��̟N�l�N��M����q6�l���^��|��2C��/�y�=R����mOԫ��4W�E��?�.�r�����.Ӝt@�sK87a�$擥�h�v��Ga_��4��|X���M-��Nb̔�9��j��>�x�V�7/�-�xQ<��X��ҹhlt�������_g4��E��x����A� �Ca�:��/WOb�Qa�p�Q�G _aS��D��)�Yi�ŵ��;%��`�w�AK/�T�ղ��|��5�ĻS�þ,^t/"�{��li����(�� |I���Z.E������.��.=��y�ѝ���w���Fߓ, :�g��50V�o��jg˽s�k�m�����$��f!�_{ ��\%�ٟ�z�uKdg��땫��k�.G�k�y���ɰ�@�Bko߾�>^��19MX�-����fￎQ����x볛��d�����&�|��_������mE"���� <�H&q��|������ӧi��N�����(XVr��l���q��E �C�2��P���^�e����L��Y�;�bK&'�-	��J�rߖw\"��[�q�W�|�8e%!Rn,��/�S]��f�e(�[l�aE5��;"��{���R�4@	��w������\饟1_
|��[ˍ>8�^� ��Y��{$��F�� Ld�����	����q	#c�K�R>��D�Z�-�PD�>�sʚN�~eF����ǎ�����Z�7�ޝ��=�櫁�Ư���8�}yǏC���� s�i�,�#?�c2�;��Jg۬9hf;D�+ .'�(�0|UZ�&�9bǷ�Yܛ�z�;y������+�wE�q}����\�F����.���\�$E����P7�.^�6���s+RB+�E(�c5�C�
�/Vg�͉L�0�����	�D�v������c�����A��f	0�5���`%;Q}7�|����l��7X}�����#�S�� R뮹F��^j▉v9����jY�S��Y��	@�������K�7nD7�P�.�YI'���AICM�қ�y���Z��h�^�Z�v{�v����i���#�]W�4�S�.D ��ɨ�b��[z�B��a��^�YNz'�f��5��.��+fu$�PO&�a�|�	���g�fL�I��g��()��#�8��Ⱥ���s�vrӖP�M�t�2�L��A�L��_�"��VjlA�f8����R5@���5�J\�L�t���Ɖ2-+5�#����rc�:��Ti�)I��c�ɋ*��D���Ev�0ڪ�5>����9��G"��GW*��5ϡ���#�jIX�$�%J"��0#�k��E�3+?:c�[��S����3pԄ_��{��լF���k!�6_\�	��_��=�l�Q?��V|y�����0A��yň�N�D>ĭ�)�.���$�Y�6l����%JY7α��ed������*���A4�:J�mU�6p��u- U��Gf����#O���-p߃������;��MT�2L�������xzBV�˰F���}5�S��KG!�I
�G�_ϑ�'&u�PR�2�z�Pv����Y�nuwy������+��D=�
'���8�i��p��tt5�6b�n[Sp�?"��N��K�X�������Qp�om�	f�.�Z���]-6��e�C�D�����p:]�g�=�ڙ���{7g-3�'s*��20D���^X��(��⼟��+FYY�}�U�7+������7�E`m0��e���Z2��'i�|�8�v��iɒ�V�n�eE�0��Ï#h�l�p�����;��c�RI��Ҥ9ė���\��gpZ�^	Tc��뻊.u�q�(}�ɟ���u<���u�Р/��IfZ���[�UaN�f�P�lJ�N�<YS!j�v֟"2$�Y2j�R�p�c���������kQw�6
�Cp�E :w|[k>�b�����C��/�1��A�jCLD��l�;��]�x�9%�[��ގ ��!057];Z����b��c>�u@�[s�Q��_��A�m<9�N/�Z��)_n�Uo,F{�� M�����<�!��,��&�[2�)�,A�%����f��d���,�%&����
)j.ގrPg�)J<�3��	P�b(�X�t��Zw!66�]�e�py��`2c�\��ج+ݎC+��rh��>��d����y�nJ�W����w�ä�Ď��Y{P�#�9P,;yiO�g꺀OB���jD����8�!�����/8 �cnvn��N�8���J|�g�?ᜃ@P���H̻Gہo���{1�?_�� ]f 0���c�ɔ!���n8}�Z�DV��5y'	��K&��t�<7��?(�to���@t��۹@��ש�N��,�o�q���Cç(�R�c�o�'�X������Ʌ����]ϱ+���=�-�96��r寔Ex��r�[,�_�����L�D��;�QCXO֏|NB��H���܆븙c�)�����D�g�.��F�}����8�"��;�M�Ŷ#����˘���X#l���v��\��4Z�F�f�u3�����Ѳ���iY�;�ؕu����i��[��Z'�7���۔�{�&�5�x������J����D���a��y�ޯtD/ʔƧެDp�jk?��"��:��2�s�-����H�^���oLU�eH ��6�zn�� k�r�����U�l�r%�Z�6B�NC��2�r{ '~�5�wwK�����
�� �1��Ć4�u1F���]Fa��RRN�O�;�
;i��8����� d�H�x�|���r�����	a�h���K	���L�ropҁh$ͩ�������F�1F��l0p�f>�d	5�;q�셏T��p=�HP>O'uA�$l���o��w��}��U���dV*��t�0Mg����J��^�`��QvZ��iV���vg�j�˂^��~�3}b�s�M�����_h��f�XE�. F��a���ֆ(��<C*u�}����c/���R�V��7���
j��	�ԪU����S]�&�Qhɐ&ƚ �Fv��K �����#6(c�f<f�U�X�Ԧ2��πN8OJ��_F_c��ZRlT�G�^���s�J��!j�����v����r��bJ����K�c��t�`7<�N����>"=���������Ǳt� }p��Du��K��?�<�гd_>�E+�P��a�#�:uC�<�� ݼ��:���
���`�ƕ ��y�<=y(��q��c�w��J=rp)Uܡ� �oE���|g멋#�nux#���Ē�~y�/wl�u=����E�%���|���܍w H��N����V�e�����/��&�D@[�tQw�T��K⤼F�rw�K��g�Ҍ��u�sI���jΦ��z?��"s8ԵC�ϫ�׉���z��ޗf�[��y�`��\�d6ܙfR�/� ;�3t�LF�����>�$�L�����Ծ��Y��M�V�ॣ� �yLj$��/�n���料�~����)�u���GW��S�3������ғ�5e�?�D��.��[�x��B�bZnEA����I��YN��Y?�!,V�i��h���lf��J �?y�5��|�WG%Og�	��[	)�C�tzY9�#��Lz�wy.�����f��@�����_���.��x/�&�
���N��F�����}Mݓ��_/�yHB�h�O�\��:(=�D%77������[���b):G�Bsn] ��1�P��)�p�{�	a�VO����'�4Ei�C�<xH�^�a��i�+�Xܢ�#�a����>��YR���K� ���"��IA`BK0��j��u��Yp՚rF	�n�J����bV��:�X�5��sC��[���r�A)d&m�1�N�pN#��ׅ�֨OT0C�@�'9y�}	����Ƭ�'y���f�XK.VTC�]�}�������k���*�*��ƽΈ�0�1I�OB�H�[nu[�
#M^Ŧ�9�-Z{2��L=rUDY���Z��!O[��~�s8VD�U�2Ž�����?�yb9[B�ޮ"�^�:��a��5�a_���c�o��V�1%�6���u'������L�%��[�ӱ�c�J�hߍ5��M[��'"�[B5ֶ���Ӫx�%#x�^β���3�}7+��X�o'X<��fA_ �JR'F@R����êtP�u(�(�����7
GDs��Ii�a�y��������쩁K���g*����S��v����Ӕ��)X`�	[��{G�OJ�sS�LQ�/N���x0^)
Je� ����z�Oʸ@��!蕁�N Fz/���y����J��\k�H��~f�'��:���b�K���)��+�����9��lKO$qݴy��:�u!���BB��@��nR�?\q�M!����h���E��C����XM�\�R���Tɐ�BW����U��{��-���_#t�IHgQk1UvtA�$�]
ݎ'�y=�>RM��������	B������[l4����@e���Yf��(tL.�AU}�><�Y�uIH�_7p�a.nMJV� �[bCA���M�owwi�0��Aۢ/v�6�}֪j[�1�W��ܳO�&[tG�,q�� [4��w�wʒ�z�b�GV�!�!o�-����߯8G��<����x�3P6^��\I�n��U>Ǽx��IM�ܥ�u����y�@I�aNv����s��� ���H��� ������b���2i���ܴ���:���m��}K�����3I�W���>�d�;Lӭ�lm{~�cpY�����U{��p�R_Zv_�������y���Y�[~Qx�	�:f��Y�
S�J�T�v�����|	�T�wo��d��5��wτ������^#ڴ��=7-[�چeK)<�
��vh��g\�>,���Ϝ"jR����|UV��'Y�O�	��L�l3D���\P�j|5ZJgi{7�h-_ ���UAi�so�T0�y.�C�f�(2Q"ֹ(��|}���YT�c���龾M�XIH��5N����F��� s��a���XJ9K����H�]:⻤��9��y�]F�:�*��L	^3p	7�Դ�ea:
���q���.�u��5F��Ǡ��w&ne���%�K���� � U���i����WOxH��To	r���I�W����B���U�zYQ95"rb�̮�LV�y�b��������yEZ��/�_����ـ���u	^Wɕ�ЇI�T�v	����?$��v � rh���`��t[�ZH4�G#�$�2�c�-���2�%�I������H���po�܋pv	���W�OQ���=6�I�d|\n��o�ZvEY��?>�t��6Lhǘw�dxW|��|��ɶJa��|���u�BƔ�d��	ZolE�Q���s�
��F�p�d}��%&p5���ڦ�]Y�e��㕴j&<��QLQd_�zQH���'	�nW��S]���^��:
�2��zB���5..��=��b��\�F�oN�
�Ċ����?Z �9��������I G��4?Q[�hw21b����4���`�P� �8kF�+ό���i�}��;�ra<W;�z,Yf��a)���ˣQ�����QnO��i�P=
�p ;�3Zԑ�ۙ��os������5G dg��1(���4�%��C?!�V0z��"�q�{�2f�V�K�ZG���9Xy.�@4����Ht2��7��;[��K,�戇,hog��B؋��!�����H�\��Upx��
����3�syK��|pA#��UԌ�%�����}����ף��T��I�"���Bj���.��9���R��q��d���J���V^b��q�Iق��FKj,�uiIR<!Ǣb���j���S�k؛��G�抦�:���o�v,���^�w5�N���3:E}���F˝_�R�aە�=�����"�uv�>g�9�%i�NT��߯@�S�{� �\�yE"8�X�����a�;�/U�o�>�g3Q�se����1�������
7�Bm��Ӟ���vt3L=0�0V���/K1�"�ȉO%�}?��[ui��[��S�����}S�s�1%'���O�0"������%f�=�yr�
��V"�8�N�$v[�km��A��������	�EN�|h����nP�W�H#y�yw4����y�X�$��]��~��m�Q���a�c���YF�T���oKM��׀��� (��H��Vn�NX�L�VdtEMƑڸr�k��6j�WF��.�h��mYh�t��qcYd������ߩ�e�0��j*o@Sx.z��KM^��'^>�ף]��#�e��bƧo��ו0��.I�#�� ����c�`.�<��U��B�i��pOW�G� �KF0Fĵy�%�?+���*q���>��\����7P���W}��p5g�TB�E�id�Rִ��=�"��z����ci\e����2��"��|o�1Hw�2�T<�M�4!���`�5&ɪDQ�<�~3�*GV7���<(���U	����{��k�4�8+�v��A��ջɼ�$ڼ2���x�LJ;>)�G��wFr�?곻��5c9?�>L|�V#�vʭIk�1�T��e�
=Ȓ�goc5�����H.D��\C��V�q�F�$t�.�Y�Z#��0w��O0�*�讜����0��ᢷ�NsW��)�6�Z5��J���J�5���z�����ⰼm�24I�o�G^�����Ո񔭃���^Թ��E2(m��@����w���h������9%�+���{�>|ڄ�v#V��XMvD�K���Ă�o�K�)C�rwz7̓8�T�z���m��[��AEX��NJ�j�e�%p�������}�;-�X��m���t���F;�[��t6�	T��rbrF�!L��"��Qol�p�7��)r���IHԔw`�(�|Λ�,�\bc�k��`�C'o#������|ຜ^��S��MT��{DʝNΰh��ў��Y��9��2�����U��aa����n6:�31��S*gE=���J�@i�A�AP.jy8=Ԡ����.y�ȣл��2�9�]�x�ន�jP5f��&� �2��G�#�w��#h님m�U_��Z�0�"����s��=J�m!��xp��u��z��o���q?��%��k2������wpɘ�ͣr��S���_��zh@-N���H2]���CK�7^��������'Aޡ��V��>!V%hQ#�)���1�F���
0������EO*T�nA��|*m�P�ܻSj�Em�'oLm-��GP�J��d��
�a/�6�
��=��EP|���h��n����x]ZB~�1%������p�
T�Ae�e�[���4��8Zm�o_�~�e��+e"�*�q��ykǡD�'�;"�@�K��Xl��͚�TsU�v!��da��F���yr'I�<�Q��?��N��	_}?�ܮ����Ϙ$M�����-u�D�`�Q��x�z�e.���RJD���ͯ�2{�g���H{��I�eC��:Kk�V��T�K����<�e�&��`��(�/͡6A�m���:��	-+U�,����[�7��zqhh&[K�(2���la��t��k�Q�&�8��
j��ca��݅�gK���F���P,q�!6/3�M5}�[ TO�����5W� ��_<))W�x���tҲ�J��!�5ݛt�Y}�&��n�s<,t`,j��Ys
Zž:7ܾ^A�Tff�`����^<����a���Kf���?.��c��(��*��.䒟���Y���D��8gn�ܷ��y����fqe��:AE����X?��G�j��l⬖�1:4^h�6Vv��b��r���CaA� % �V�M͟Oi�T[h�z�jz��［-����MS�=�(�6�q��wÃ���ՂX��VG$�{��~P�s,��5�5�2VT�� I�E�ab���C��� +�Y]iR�sh�jY�E ��+Mg��]xA|"n�r<�\��鮍d�-�/gDŉf~e�}wH�ۜY��2�17�V��j���Fp�Q�=l�)f9�S����Y<f�Z��xJ>��[>~�=L��K�����Z]g�OoVɃ)}���˕@4�����X�7i�!Ա�1DM���O�x��Z�<�:1�E�K��[�%����ѓa�=;�N�	h��mm�ڂ�)��F83�]ؚ��2���b��uy�<[rg��J�������n_�z�@����@��Y%#�"y�mm��������;?5;�|;�%_�U�U�+��2���Jb���n�7d7#����)7����k�JMo�z�L��*nA��	qbpA*��rE�1h���C�v;�w�K ,������=���	e'L�����{�%�(�u�9�-���&^��!qDs�C��5�7�.N�.��.���RD�M+�l�87�7�Ƚ"���������X��~��hG"Tx!��?�0e	�`w�p�8k�z��d���Q����E�t��`�x�|e[��L���K�zg	�����5m�j��B�?��g����͸f���&��_{}��.ࡴ��ŲU�����t��]���*�P?:� )���ۤ�*�es*V	��,�+1$��Ӑ�Ѣ����-]qbT%����T����n�̊0�W�ϱ1�dB�h����|�_b������mu�JL\�z��?%y�n���*�a6O��Q��M?�� B(6>YLq��]�Y��#6gS���ei��.A��]�t��S�p�P�Q!���e���41F=�k�/[>�u$ޒ}�^sZ]l(�����N�H�c��B�J�P�e�%J|~nQ!���x��ŭ)Vz�Z�4Y$Z�����LE3�a�nk��uK�v��v�|�Wo9H<Iᚸ��L�`�?���kS%��-=88^8o���6��8H��
���;d�5$x��
0S5'�8�RQ��em�W&� ��wL�}}�8��߱�B��-�Go�`����+i{�MԀj���ipf�C�jŖ�����x?'�
+�O�l�5�~F���n�M@K`�~*a�ɫ�>���*�c�����>�I\�)��x,a���#�BH��z�r&R#%�Muн��h�^�m"��k�a��{�L�>/���B�WC� �E���e�o���%GC�F�-������"R��)W@�B�&8��Q�~ǝ�5}
�a�J�'�a�$���2��)�1V�w$�X�rC� ��~Q�\|6G��׽ MSSM�(�{5���g�Yk֜��u[��H��G���Qs��b�B�}�)DAm�Ũo�.gBZ��o��3��f�j�����y�^���"�Eň��1H�G�t���M�&l�;2A�����,}�abg>�m��r��������d����}��`a�]�]�EO3�8����%`I4vpj��'w䝟?'��04�k��rt�yaw�	�_ؤm� oV��4�G]��B�²�n:`�E(�_jF�r�;�f���ƇE�� /���`HD��@�o_/[���#@TY�>P�M��Y[a�o4��·�@��P2jR3�<6����!G�\(H���D~�t��/<�������(z,v�~�����J��{;�ؼ��%��ծT�7ٚ��CƴTv���[�x�$�6SMgڅO�
�=���<K�V_���;8�$r���C9�yL}A?"�M#PÊ ׁ�/m��${��\/��0��H�{Z�6}�\/�U�!�d"��L�՘�o��{%�{����j��
ւ����uD��L.�TS��)=��Ui#��W9�L��pm,w䠽�G��$�Σ��i�c	sm�2Aq��?[I��yJ�b|v����[�=�e~;��t���=_�r! �P�g�ج�iӝ�����=4�$jp30��0)�����B���6�k.m�|Iwq�pflVk@p�D��X�G��1{�����]>��/�qy�l:�@1���N�>i+�q�p�9�a�&G�=(�_/�SI�u$�׾�8JY����k�Vj��:�� ħ�s��dVRb��34�ǫ�_���o�e�X1�����V���K_��F�{G�j�&KX4Su�|�k�$�����b�e�H�=�1O���R$L�gi;wr�M��3�*$ҳR��Pe6<G�^tn�����Ug��)�c�O��a��dЩ�~sY���	ȱF/7�Kugv�%�} A�ۮ)o��y�n���ú�&��-��^��߿8�YTU��0Vz�"�����\4樻��+4�]�+��"�j��T|��H�t�1�i�A&�m%4~X
�5��I�Z�ʮɦR�*�?ΰ/���YynsCWQ��B����;b�Y`���z$3�������ah/�*Jk���՞Z&Z���L�j��AZ����bS�����b��jyr˛k�M�L����ǉ�k~�����G��j-����z���)x�P�j�)�iK[`4���;�y���L���2>��[���۲H����C{��0ss������ ��S+$vv�uv��C�]Xn��F�1��}��R%8�X�7����e.~^�/�ؗ"�m�� p��']�I�@![�0��9(A�C��}�?a3�gy��҅�	n�	O�`���9���xԞ���_Tw4�����M��P����a�(%d,�)5�V
�
$U�Z�a�o�u)@o���7L�G ǜ\6|�
IL8�w�vh�S[���F���
7@�{������v.����0_5����T�*�&�&?�Z�g�4ϟ������ɻ䉲��IǨ��-j�ǳ� Z�&cC8�	�f�r�R?Y����3��Mtc"d��,����䁦�e�LAf��i ץ�vS�����=��"�`���

�mx���?|\_
�r�������M��Q��F�j��nۼn,'�"�
�0*�ȏ�x������f6�T��;�
��yw���uP��ɏ�N�A�3�v���`D2�D|�O�E�D�3�YJ�`�t�&I��q�̫WYM\ʙ఑�c+�O
bݼ�Δm�@���n���e@Y��Wi�飥zn ����Jʈ�#ˆ�Ԃ/?eB~(���t/J�l�o[9 #<o�}:;��_�:5�>Re�>$�>�q����e��яq�Z[ӡ[�+ݣ��xW��%?�+q�>�M�3��{�WW�����DP��г�P��o�E��DFN=��3�e���|��ʂ�����u����^�jnP���6#T:�>Hb���o)����k�~3h���Jݓ��w=W2d�����QB;"#��� ɢ5	E�H�-�H���Đ5����`oLBo��3V"ނ�4���}��[|0]���zǕ5�� SY�s�Dr;�� _�E�_��i/m�_0��6�A��㷚�F#�!����#���m'  ��,��~��$*�݌۪l�0}�i}%������9�	��(M%�����ەLo���HL���B���A������:��C�����^��I��y���%e2<4,�ҊX��H�ܛȼ�J�-��<(�CN��xw�>����%.}��6Yt�6&�H3}�Χ���G5���fIW�-��$;}�+j�{�e��J[E�+{]�_���#��œ� �K����2s(���.r�c�'���7N�9�-X�`p���%���^��Yz5�6\}� +�ΜX�>3� ?��j}];\�3wvoY������uB��j��1�/dw��g���V��#i�LV4�B����~l��/d%� (eO�au�1�����C	1sR(�u�2����01�UB 	�iu_���A�ɩ�T�Olդn�5���Uʋ�ٽr��JY�fzW���B6�W�����7h9!c�}��-�64mZ��@\��pz^J���zW���^3�}�������"�ud�P�:'b�p�.e�sg�"��0��c���z��?�;��#R/��^�{r�:�$�a���~�+˺@�C_�I�%���I��kz­K��t�Z�d$�Hj}�LN����1�U��.>�`�;�q���d
-�_)�	�Pi�ƀq�u�X�4��b�����6��:��v��/�G��P���d%͡��l��}��U$��ț6%�c�T5z&zq@,%r���g�㳆oi�L||�){�(���M�tֿL�q�A�1��qAѸ Ki�Q��߄h���0rn����6i��_�����EY�vH�
���
?�V,E=�OW��wv.%aZ��X~T�k�?���-��VsV�K.J΁�i�a��L0Q�3���.�`�rk�� ���y���l,�2��&i�\ήv�z� �8��=}�5ox̋������͜�mK��E��^���i�֙���N%��I�kH9 	�`ε�#ޜ�z���/�n��[u����L�x�g pv� �9BB��w<�)/��3`J̘Ɖ��L<���5��S�:{�{�ݩ�Ő�e�WJ�{�bC�����LG���b1k��ʀ�ڊ�$�̝��T��@\�$ h�'D�v�ࣶ��������!�¡���E��r���١x�����)�k.<�[��i\�"sa2��Z�>F���qu��ntQG�.9kK����m�voٯ��cK�ֈ [�1R�� �MIp�5�b3�
�<�
q=_�O��@��aͮ�
A�A�~��@�������֤�JiXY��9=����W	���).@�UE��b���S�9zNr^գ�"F৕K�̷sM�;���Ue �Ч�"ݭ��f������� ����m�ڣY��kƓ�����%��)�J��m-i9��#II�|,U���G�US�c�}D�J&sa���_5�NV���V��؅D�ҽ�����U��k�Qh��Ƒ�$��|��Sr��i�r�E!38Ce�D��i������s,�^L���kW���q��I'�p��Q>��
�U������!�&;=bלK�������V�#�
�-�Ϙq�e�0A�8{*�ۜ�7t%13zث)�,� �'\y��{����u�h��� r�����>�`~����1��p�S���!�Cg�u��N���s������_�F�ޮB>*�J.R �;Io��� �[��'`�P{0.���e��)"��}C�0���?���Ц����{��ʨ���>�r�a&���՘ R�u�~7� �*�xC�e�WAn�?4 e�+���97��]�3�+�W�G�:��8B ���Č-CWw|����-�.ڰ��ʧ��1]�6}��1�E�g�}�h�WD��MYQ:� 9�N'�bE�u �s,�ƙQ�r��"������{^P
��e/�����h�����Hz͝3Q��tc���4fB��[_���C�V��}��Ť"�c ���=�t������͸�S��?��J�3�X�!H�&��b�M"ʂYڇYq��6��|<���/?��C+�XX�u-��r�0ϕ��J
7���_߃��C}n���f�o���V.�{�!�}e��~� D/7(Ⴈ(F�J���yey��z�o��ni<��y�(�ّ<ы�б�_������:��������c����}��p	1�Zb�\�=�����:I�u�%�� 8-�0���tτNe�v�=�5��țW͙w��#ű���,>��Z9��s���"B��p6��v9=�� �E�\:�f.Yl=��z�p��ٟٝ�\��s�
�g�x1Ztz��jC���~����{xA�11��$5��[`{��,�Ԅ�+��lU������C-,F&?rB��y�2G�)�3]E-e.Y�]fњ��o^o%t���4n�Ԝ:��M�4��Z���	���P��]�0̎�L�`+R�����NH�f�-*�>f0���n���A@�R��4�3����*)g�=�Z;�\n�B��*�6I
#dH����"��spH��	}��D�K�u�W��vG��N3�Qۨ�
�)��VM y��
d��3H5�E�3���՜����)ݟu����x�@��� u��"�p=���d_�qں{(�y\��g�1�2�����{T r+�kܲ�G���K'���H{&x��)�x�N?C�u��Q��Q~W���[�|�����c�'�
��I	;
L�
�ʁmb�qZ�NM�;��b�T-i`&!B�)��30*x{�qs�,RL��! 6~Q��M� ��(8�����C��^\U�~�[�+�����hZGQm��u��𥺰.>"0�	i]Ԭ��A�-��4��"�m@�6��x�"%?>�n�AózȎ+O��=v����	�&U7����@I��z?�� |?��p�=<OPI�_;�Ucԅ0�tt��|hk���9r�v��?�3��+JD(Bd�p���IvZ�(ּ�_����"�[I��|��G��f(*�)��u��鼤���#S3����nF�����ۥ�(���5��]T����^~�[S"8o��c�6�����X��8�#}�4�];��O��݃M���"��6 h��\����u d���/��=�kC���tMӤ�q��2�P+y��&�{�y�������V��~�jwD}�tb����)�������ŋ9���H2�BV/DM�fy:4tb\?Qթ�Z�~�������}�*��^)��~U���=+�"��u����?R�\��9��ֹ�/�A�{7�.m���-�5����������R�+Z�m� ���O�Ԑ�D�2����<�ڬd'�|Rэ6W�Kf�爗pU�b�S<�#���j5��?�׋��u�*��/�o�*�.�oB��b,�n�8V��`WU��0k�k�m�ᣢdfc�b���|++g� zR8Ŧ�D}��	ۥ!(و�a��p$��p:��OTϑ`7l��+ G��i���H����B8���>+��"#c����f�_5�8�7 �>�L�EI7��ݎKi'��`�3G��k�<FWmç�o<�g�3���)����߿Jg9����Zx62�mh��?�p[�Q��1��Ќ���i�UWچ?�6��D�� �iA|X�{�8�$�ô���=IV�Q3<,�11��e���Z"�����v֣υJ��h�
�`qş�*(xZ�$�����g�zJ�ý���gaS�,�Om�+�¼C�M�d<��AU�;�u�.[6�8��mܶ?/{�ٯ�k�u�rl�J<��X�C[t$�
$@v��FL�X�懲U�+I�S�g���4�|,�EG=�q�;D�_9{�8�����y�ү��|_�g�ZE[�S$�&�".��-�F�Cv��G��Hrm�ĈW�f@�`�����*BC$�f��K��p�c<!S�Z����+�0k��"Tr6H{�K!�֕����ڼd僧���?ς���>�����?��:\t�-%FĦ&uJ^k����+q_?Q��E���鞴;���yg���IV��X��������z �믅v��d)�{�ȏ�^�����&n�+�E������ U���$`�٠�L��m`tg��ݿ��������{��=�ǈ;0��O�Y<���X��=�Φ�Jb����,ٮ�_�%z/����QO�Y�V�쏸lʭ�>�x�,��]Ιh}�����$-z���7��]����qh@isF�x߹9j=�S�XI���G�� �'�V�z�DI(��[:ި�e�S�o��Ԃ-���o�Qr��e:�{!�o�3m�|���2"�ζ�~YaZ�K�y�W� z������S����XŔ���$$M�==!�H�G������Sʀ���6�@1_��.��?��5@q�?�ة�.��-����hֻ1�>��'ȝ������;���B4x�8zw�~�����lkca�Ӧ�[��9#�r�pW| b�Z�(P ��j�l�x�lʕ��n�������b�8�=�	�(��5=L����g��+tQt0ϥ��iv�|�`�� ���܂����l���.��fAC>��?�)�5��}�^�>�'�<QO�.<��-�|�=;�ШQ�n\��j�v9�xF�W�8�U�ߦ�|�ӔZ:�7���������\�[�>4���ۄ/y���q���$[��#I�8n��4xjkv&x��e�����Fx�/����gZ�/?�W��.����h�]��U]�X>J�y�ti?y����LJgS��E�;��y�����|g�72�hl���Z����M'+!�C+ý/E��Y/'�ٮ���|쳏��Xm��{#l�%�{lmУr
1jc^����.�As�	�JD7������+�5�1�찭�ԧ�w��y6�2��Y��uw���̑/�x��u����vxC�`�Ik;����K�/���E���pI�	Nܨ�<��㢝��V����5��h���P02�^�̵���-���4����x���`8㙞�mk"(��'��L�j�pRPƧ�������]�3®��Nn^�Z�)`p&�kw�����h�������,��6�\��x\���Q��5��O����?�T�X�������� '�j��z+��4JAT�;��̺F@���\OPqV������E�0���I���z���4�߸&�:+���OP�Cg��`���'c�L�F�f��c��&��ňTjԙ�M��yZZ\�S�3@�%�)h��a��z/��|k�Q����@=��~��4��ru�#���_������<KO��GNB��G%�����Q�[0�,�F���W�����,s ���G-�i_D�D5������-�6-;�81LOր�(��"�g���{�+o�&�ͨثh|������lk��p��k�'Y�ɛ����fϳU~*赻t|&+OH�#+w�yQ�=��B�HQ�M�0�~��·�\��]�m6��i��6�CY'�?ҿ��RnO�PӾ�r��\~�d���82|�&D}y���n1)��p�r�ea7��}߂!�u�����r�*$�Yu���y�5�����Y��JHv���Y�S]�iX-Z�K\�)Ř�?M[���=���O�G�E�q8��Ϗ�as�����ㄽ-���s�Q��r�`�FK��h�0F&�ð'N�;R��1nK�@�y-Rq�A���9<%�B�����2�=rB�p4S��
����)Z�^9h�vj"���@ME�q�1��O�,���ãc�>����+Ӏ4�o������C]Y��4H̾�������`�C	GB�I������!/���
��@��no����$�Ւ���K�MJm^`���ܙ��}J�|�q�{5,�?`�i��Av�@ߑ�d�5��j��at�����%Ďu5��Һr%9�{�c(E�J�%w�ժB�|��6�I߄c3����xk{�f�]p�_Z�4$��٣f%t����\�����p�y��/��z��/-q.@�i�q֐-�<���V����i�Ʃ�ַ�%i�Ȩ��F���P��[�d���,�!Z�~���b����ǁQɟ{�}؍�����;j�tO�G�� ��6� m�E�f`�@��?LbT�2FF��R,ݑ���Y���������5�8d��t
pk���*�6��J|��oK/�lƦOX;ב�K��͡�0([�s���-��s�!�gg��������R�ei�;���B0�^��Q�T1^,��:S:��/�����ss�Q�į bȕ<������Ć��g5�К��!�V�N�����}�C�Pm�ՙ��!/M�+� l�T+�x+`�fp��~��P��YyR�9�[½d�K��ḭ̆Ih�1���bR�{��q��IF�z�`@��!�>�t�/�Ŧ�^����K���)����M	��d�ߤ��í�I���%����.����) �+V
T�oL�f��(&d_;�\6�;�%'����L8��;x����a%��	���N��gk��/�#8�u5C:��h_�O��1���k@-��������ʋb�#�LE q$(�_�ͬ9� ��X��_���I����B��od�~�.��&~;�f;�/3�PgF�$3l���G����{Sڎ�����������o�^��������e��s5������ػ�?�8K8��CY_V3�����u��$EN�٭�������� ��t���%�樂Đ)�*�UVА]���eoS���R\�ޅ�r��HY=i,���Z�ɘ�8+Ј��vֱk��rw�q{���b�ܽ��١ꦄ���r�`K+p7C�D�s�,��&�����t���s��݀o�Vžꇥ��"uY������e�8u��5��y��C����0t@M%��Av�?�%*m�{�J���2e$�Ydtғ"�<"6gÔE`�����^� �����>� ���\��z��,{K�)�fIb\��^8��ŵ�Ւ���gq�07�gjyd����$J�R�n�\��h�7Uu�35_��I��?F3�Aگ�T�"�dx����2ː>F��{�w�=��v��Z��rH7�T$�w�T���4��Z{<a��ڂ^��ڛ^��0\�8�9�p�jѲio�:N��d����/�[�/E(I��9�Ȉ����-�ZPb�o�Ũ���XA���]�j�.�Y�4�3KmEE#�1�b��E�I.�!�h� S�s�7ˉG�6x�C�~�zػ��j��\K<�m섏j�(�$���4���K����(1���������к��JE��Q���e~h����<�G��nK�"�D�aiW�f��!>������5�T��'���db:@�%V������=S10�έ��(�mz_�^�2]_�1������i��Ác��D���XK�;MT����%���:wQ��8��'?�Fl"��'��ʸ���k�L�6&�"�#P�G��S��`���h��,C��jv��1XR�'Iтp�I��D�� �q�#Qm4�.��o��pj ���.ym�N��� �+�&�W�,/���N	��ugO�*��ZE�yI��t��"h�;ak:��;KNއ}�V����ҋ1���|�0%��2}�+�����)<j�9`ѿH"̵���cpO�Im��a��kD����g��:��]����=�[��C�,/N�{�o�ְ�[#�[	��/�c5v����B+���$Z�Vű�����)&:^�/z��Ж$;z��)��`8���9�g�h���#���B u�����y�<�H�xa�׶��
�^���>�c�g�����K�����?�=9��E��h��6�e4u��#YG���{��[��OO�a���O����%���j��Ғ|����7��)�٦<曙�0�=\6�Xa[��߳�������:�F3�G�w!�����"މ!�qF�S��AzK��w����iI{eт ����\'�o	���D��@��F48.��i��CEV�[���lɓ�q��PI�PK>0�Տ���o��c%x��e�a��"n�ʂ>����5+���Oi���BA��փ!u��I����
��M�]��k���0QD'����+�q�e�s�?΀H��4��=�z;혇�2<R����+�qDg���~���v���(?K�%�[�=�U���������=���ά��X ��z}������.�W�C���B�r�ts��́R�:��A��J*y�eҟ��U��V9eS�$l��nPi�V��wo����M�e��+]�(�Y�0M�	N�c��ؓK+R�D�*�e������Z#�����@S�T"��,ֈ��gB��������!��dT��1�|����K8�>u�4����gIL�%삚/I3z���CN��|؝�>��Ӂ�j;�#�xˀ���Q�E�۞-���IeA�Яg̝6�GAS:�ȇ��9���drO1�C�~�jn&�M�� ����C4%�X��2�3�Kuݏ�a��_�J��/��exJ�M��(L�E�>J�����d����*��ʞ�I���=<ԏ?��R����&���t�pv,b��>1�r��^�N����Y�b�t�Z���@���	0Ut�V����-&$�pD�� ���ս�ݐS8�te8.��%c���l��J�>���{���#fW�ʮ����`pBk����W�0���P�$�[�/P#����Z���Z�jn�N�W�}^��yI]�W�+G'��0�]\�?���|���v���WE�ZH�y<����f��}q�D<��'8�{RѻR��|��<�Zaל����a�e��+s�G�C*� �{m	u����<�R�׋GPʸ����cr�u|sWV��O�L� ;x�Q��m�v��=�O(-����wY9��f�C���#�}�~���Et���P���R�wii踟�5�_�9Fo�Wq�ٽ�#�[����Ƿ��T���h�@��_)��f�J}ة���W8_���5j���W�QX~�1�K]�cLH�xx�rAJ0Pz�#�r�q~����f].�iC�7�P<߹���$��r��4;ň[�|�s����/�����}�=<@�l��zh�n7=U��v]����&��s�,F3^�+���{�ћ\�Bh�R�x.d !� *!޾y�֮�=IZ��v�!�/H�ej7�y˜�LS����=}]��̗.R!������6�(T��s�s�R��L��	
�o��'�g�[�Ri�RΎf���`iJ;� dT�|��)���:�߷�8
^��j�}�Ĥ��EYB=e�'k���#�z��|{ro�|���Xh�@U�E�����>�|DML1i릏,�M8��~i��c�g� Oor*���PrXe�N.>]^��c"�'�z�;��]zeQ`�=��~˄�����"/P0����K�9��-aǔ�8VI��>���Z��x��8�%�_����>�)٧�m��ľHB5��l��vޠ�<�I����`<l�~3��a ����{�x��η��hs��9V �(�C�?�z&qv���|�n擿���2f������e>�A8!M�9&�(��́��|��o��O�V�e`����8)G&p
P�N��&���y�Tש(�<��k�W�$�2% �)��hȍk��="�A�װ}��� ��wy�:���yJ����� ��hB�F�~�iS���$�%A�<�P�gٴ����*��X�W��^u��~�8�D������ί����}��:��4u�F%=�bO�����4�� �i��k���.��pa�N�����^���U/V�j	Z-}�<�����`�u-��2��]�팃���M\+ud�4nE��W�Q��?5��)�4��}��b��4�G���'h�P��/�%��~9�)��$\�#��G4�}	��<���E�L� �]�=�лu���r��(�M���`�@��+Bʨ�b�ɞ �߆����5y	�QLG��|su����B�]�*X)�7@�O7��C�Ȟ�Ăz��=X�1���!�N�{���_}&ԇ�H��H oD{�u�/��:o�xuYq}o2ǃG!���Z�@�#�xjg���ږ.S�Ά"]�b���ϼ�[�t��Åf����8���l-��hYMCөQ�&c��O��$l�k[��c���<e����VQ_FŏB�Q.�K���<��A2)��j\v�/�:�f�w%�n9JYXX��O��Cto�_�+��C�
+�䇽R�zٙV���DA���v�=����6'ݬ.bq��� ���VE�R�>x-IyipP@�8T)C]�[�g�c�>�a�d֒��o�k����/IV��D��:�\pkJ
�@e�G,��O��0����F�o��v��>I�K;��8�d��>bi���b��$�~X����n^zh�(�B�^�m�
/�����<w�M�?`���jJWg���o�Z���o���'���~�Q��I]��&��?QT����"�#����ſU�+���s|&����s�t11� �u� k=����K�99���u(�f��H��Q�.�'�P�̑w�5W�ba�&�v���0��b� �聾�=����{L��|u�R��,���HU1��͚��x�
����n���`�,��8�(M$?eޭ���z{	��KWn���%IG$�w뤒��uI��	���6q8�;�~d9a������/�	��b�k�Q�W��`�	uq��JG�P�2�Kw@_xL��^����f���������f�K�Q��������6�8�u}���$9$��EC�7FU~m�mN�^Z�p2���1�{+қ��5A�sJ"lq7:�X��#1	��I�f$K�*1UgN�G,o�Y�G�����8d:��pdp��H?I	�W�C;_y�9_��\-�P!/���2��#qyZ��@r�=������'}��1nЇ��g�|T��|J��c7�L��)��^$�Ŕ����-\;/0x���Ny�r(s������`��3G&�j��%aZ-���h�p���`K��XQ����4�-��Ïb�>2��e-R�p��++�LLbN���*/�c.���)hX�{���G��,���'��A�:*k8�%�k�Ү6QeO�4aD��>��j��ѩ�#��,�g�a�q��I�;�DL��=����K%_����d��_7�(����H�A4��x�V[F���q�ׅg[| ������;x���u$�F��f�¯�H�\�+��g��Vط;b�O{C�Z��%���|j^�o�j䥄p	,�p�qO�b,c (&f�y�唍������sumJ�x�?�SG|�=8��o���W�<�Q��I^��T�g�x��)�ܱ�1��|� ��~�\��Y}���q�gu�/�p�jV��+5�^��ڽ���.��D��y���q%�aN�&�izጸ2Զ&
 �΋��W��"����z�-)(��m�3R[.��
BD�g�����u�᭍:�K�s���?.�jwǀ�K3��b�ߛY���}ҦY�Ң(텈�1~]�ڧ�_��y�2����5v'��Ԫ��=�*3��>h� +��
�eۯ2�m�S��j*h<ƺ5*��Wi־�I���P���Ю��4�k�v4���XXi�*jqӬ3u��/�Fz�s�S���}SC����L�����NG=I�C���R�0|^���{��Y5m���5���]��ƞ� ����G���jD丏�R[�L���
�uKT��������潾�l���j_�7NV�ZX��C���K��\
�Ru%��sF�%����|"�#�?��똺����v��]�j���"Ǒ����3��x��j#3�l*O��m/uZ��π*��@�h�	w�+�V�$'�A��w��%�pcr��r�e��R�t�ͷ̙�fO]�L'�/�H��Y���x!j1 �F��^v�`�������+�6�|dC�BI��k�����qOʙ8�r-��3�w�?ް�uQ��C�'���m�����ӓ<{�H3��e��%I�R?� 3�m�945S��&���M7P�����p�	8b1
�qB4���#�R�$��*e�3�)v�w�ة&����`�x���p�Q5yDך��W�gK��nz�K�0w�_ځBNRP�A���*?3SqƄ��r�:�y0�=�mS�͵�Q�M|@���J���J�q����\#���*��Z�����=#�1©qa&Dw>iZ ��D�w�����a��3�B�
����_�����U�0�
a�m@\� dR��*�AZ������<��d%��56҉��;�ط�W ��B��}h��Ш��%#�[�DGqg�44S������#�˙w��Gq5��T]��<�WjNH��ﲚ��s�'F����Z��=A.EMb2��`o��G|�J��Hƽw��pu�x�Nu��V��a����oa�4�0�Z1lf6�(2,U�
�x�D�x��
٣4a�po�~�j��;6�֬�y�O�iǻ���;ow�$*��H4U�����L��e]���?���������#�f�T��Kn�u��Y�ģ]${���hׂ5OkrO^#1����b|@U�RI�5�/�IrbɆ�1��	?� H�*W��_�����������o!���`��{A����m�Z�_���1��(�i�xs��'����H���g4ˣ�c���{�Qb3�P��vra��d7��MN��Daa����vV޵���#�nL�����01�����x�X����r��Em�[L��?�5a�����׏�{o�%���ь-3�*�TZ�ko}�4�&g�$X�v���O�G�=nՃ�c�yԸ�Sz�w@����<���}��s�*�1a׌ԽC��Y?]��	�-9j�7<����A]0���9aC8w]<�c�&~��k�4���/>�9�����-�y]٧W K�',�~�UL'�(��f����ޫ9����V����e0���Ƽ����d۴N?��q�)Y�ߑ���������LL�U�u����
�dM��Y.in_]p5gb���s�e<�C��7���m��1˟롿�;GT��f����y�Xh됱��ɀ��h���]�PT�9�pbU.&S���Xw�����fql�f��� ��]�Ǹ�n{plt#i��:͕޴�(��L���~���k�X}	��e�4K����~x�ۖ��8@�]3���'̶6_��VH���ӗ��Ȱ��W��d��C�6���0*���F��0����;�Z��z�Q��!P;@�0�~!)�b�h�o/M��se���-�J�����'-<��*9�Y��.��G7�'�>)�jp�8��gy�o�dGY�R�i�`��bՀv��2�0v'��Q']̑�Z���lV�/�9<�JSmY�_]7�}���R�l _��J>�(&�7�j�xy~��.�$��f�y8c�s��4C�:'����M��qݨ��ɫ�o1\�6�(��7��N|��9�×��=�L}�W�hьI%���ky���p���W~�F���/�Q0����9�!(���}����Z������� �&�2xH��'��m} �'Ɨ���ꅰ�<��Q�#IU��s���"`�	�����{_i�k$���]��p��WU<��AhzO��Z��l�.i����ڜtZ�v�� s��x�$��?B3�&�, N���4�(����6�5�ѷΨ��q�=���:��C��\w��4��-���p�$�
���y�?��m��`�9V\�n��i���uj`S�>c�yFY�K��Օ�i� ͓������.[c9���R�o��$��~��F\�Go�x��G���q����w�.y���;���>�cgb��K�Z���#n�@>�%u�mHs[�L�7Y��X���g>U�5G7Q�j�r��Ky�{����_�vV�So�V�s���s�U���IU�,77������+�6��I�/�V�`/��c�ZB�W�o��؆�|��s\��6�����K"'�Ü˴ő�ֈ�"[2�0T���ާ-JZg�Ӧ����.�#��\��T53msLAQ%�O��d�����~�Br�|��R]�~����S�z[GQ� �p����4�u���D��7έ�ZX�����d�855�~������(;�#j��ŜХ�:K ..=?hsA�T�+wre7��k+]FL�p=&"Hx�z�/,E�q���P)�s��-=��@�t^{���S*[��+x��E�X7�P���Z��$�k��}��H��p���]��U����\���oZQR+a��

F@����T��_��g�U=�@82�@��^���jpr�dYx��m{zg碏��덼U�|������� cIʈ�@K��ʹnLr���Aԧ�і:���MqP�c�yo�!:�.�D��7�ぽM5z}O��_�ٓdJ�6��$w$bָ[�1E" ���AF����N�m���C`��W�*mHM��P?��T�#�O��%Es{�]iF��z�?c�$f�����zS��$S�̄�~y�����J�K��+ޙ�Ǳ�]pm�?�H7I���i��t�����Y�Kq)�m��D��>6�uE�B�`:#򡚔l�d���d-�����+�Z=��2������Rki�s�ؽ��Y��d�̝����ĝ��cS* 1�n��Iv�C�j����t_�&�����l'ߣ�ŌHG�o��i{ ��{�#T~�B8�h���5?��_O��LP���7���	\�ı6��Mb�5��n���j�'�!-9�.�R�פqK}�9�B���,���U���^�-�S�d�'3�A�:�T���n�~�(ە�1J����<�h�U�V�@��i�G�gw�ʕn ��.�|�f�'d�>P�c���^v�s�>AS��y��W��}B;:+b���:g>���:���n%��j7��"����x;��$~?���Fo�n�TsdՄ�)EE���}�,^砐�>9�=S��f<ض_��ʮʙb�]xӸ�0�7�K#��tu}��Ko?��9��:���P�wJF^�ȭ��	q���Ǌ�)v�@��,�}2w̞�D��U07&j��vQx�󘝚�	Q�rsl�Dhi�1��Oxt6���.e'�J��F:Uȋ��F��&�E�W�W@[L��P9�%hF�S$Q��/�1�嘠<"�����͕7y������{�2l�ts�|Z�b�^�N�C� ��^��@+iO���M����&���aB�(D����=kze��'`�3���עy����@}�G�n��o��SN��p²�*�<23�6�
Ṯv��y�ő���t2V�����Q��>�0	5qT�
��y&l�4e���Iʣ��Ï2FR���ےuJ`c]ICI|ʬ�Q$J�G�!�Ί����� E{�1��v9�p��4/����dC�H���"� 5<����}��S+��\li�H��D��V�9X<9(�Ȋ�pӈx����a�ǹ���r���:G@�_FPZدP��n�.ڍW����K��G�;|�i^�Et�S���lv�;H�D�ʯ����6��]S (�?y��F#)��M$��B5S����]х�{�c�y�W�=�P��ht�'�s���C�8�4	�W�����2j�zڌKV,���-�c�,��H2���r��5+�.�K�ּ��Gi��/x.�(�+��F��f�7.3/����"9�if��/�ü�g�o<�f�qB�q�m��qu�c�M�� @�0p�]��wR�%���2ˀO3kRq/(�ϋD��g����c/%�<��t�!ַp���˸�4�"d��� Zb_�
�����k���%�a�����?M���Vs�ߗg��"vZ��S#��"�����Z}<:	��	��C��9��%��n�v;�E��5� [��MO�ї&׍E%8�%a-lJ�i�@ZM�c�.%,h� ��'��}s���R&�a#�5	�XUu5���b�A�A ��	LZB3�"�G�E]
�� 9��{�%���-��r�[�o�_��i�S<���~l�剤
�����*5�D�\$	vW ��ʪY8=�����Jض�xַKT�	X)+�&i��(v��Y�9���:2*l0P����Ax� ב���K�g��c�ѣ%d�NG���&[�VΙ�`���:����.�3}��`�� Z� s3��K{�=�a�V`x���%�w�Ȍ��踨bx	���ZBiL�����/�vy��Lz�������ηg������+p�U�ch�6�Z��S�1�OS�����]�'���e���!�`q|�:�	�^�(5�(!�������⥑���:[k�n�1����429���dSbB��&D�Gԭ��YJ+�.>Ga���;jL����&G�_8E����� ��s2[�6����n�)�1��MYK.�&W�Ȏ�(u0n?sd���Su#���^Uʟ�/�b�������+���*�P���ԗ���'[��I�M�nD��r�
�m���iG�)���A�Eo <��-����6��*o� ~�s�����X�f��[���P���_@veF��H~��(pD��ַ��Q�R���Hn�
8�գH��v�!5��_���Y9�7�PlS�����w�7X/��8��=��_��U��}��&�����������)�g�V�b����Y�Hy$�����¦ @�K~<�����+�{���6j)�_P�R���Jt0�P.	Bu�\m��٘������g����+�O�/�q��q��TV�k��=q��&3Qh���+�X$��Ě��l�����$
+r� 5�f˱!��-/(G�<�5Ô�"uZu������"����=���a'DM�)�̎��ܙ��r�Z4�
lD�)2��\D&�@��bs�83��k��ы��M��^'��	y�.��<Ԩ]��4n��q��q�|ox�:��v�k9�vJ���Z$�=U�='G�Jdh9��M����D�Bd���B?ȱ\_�5Vl�H��-z�L(�X��s�L�f�"bo��m?�98-
��%�����.e��\ף��pR���R"��U�2eyWc�h��u��CC���^��2>Ĕ��F,<s���	>� ���Y�	�*?8��CA����!b�A5��7X󻝾�!�"��f�A(�i��)�[������-!� �TEΏ^H��{PA|}��0��/a��e9<�6R7v��6 ��sL��y����bj-����1*܀y>��2�$���2��9��K��*�Z�h�)9�-=q	a�l3J,̰b�$p`�!�x����=N�����ަ��I._��u��1�/�m�&d��S���0��b,��������s�+�Q���R���k>�"{9�p�7Ka=�6qغ��B��C2��l.,������j�ۯ�ś5�\�W�O�����
�T�	Ƽ:&-��P�'@�8���pDM�N�x3*�)�b�=���в2����#{�.#|W��|��2d)�3����.�����ʕ����,�M�^��n�G���|��_�l�[\����QơM�-�qd��h�������P�ū��D����%����f�s$�܅����@��H>����V���K���VN�-����/��>�e��iJeD|��Ʃv���Ǯ�sh�yM��A���tVcryDmAO�L�\�
ܒQ�+���V�>��6ם����OFǺ�Lw΃A���C��TP;�&��;�-4_�UOw��C�zظ=���3�,/�����Ф"�m*��ح���^���8���C5�	��������:M?��/��o��3@�no1�.7�qw�]l�50G����]�1_~|���0q�����{���Z��K�@c>���uu(��q3���&�,������(򘳥��N�>�]%�4 A�a�!�n�ܘ0y��)K�t��o��qe�@��������)ޚ�����MF�*���m����zmo��1�9~!Hz�����w,��E.��{�in�ؙD�;��`r��JP]���wiw��I��{J.�l�R�|�Ư��L_
��wI��_�O�ƘC���cA�ܼ!�ަ��크�P�_���CzшD�StB|Y��Y��<����E� �YȨ.�P��n��=����M�%��F�u������Xx�.J?�ojp2.�b���p	��EW�t�y�5t��iqV=���G�:=�(�N�
��g��f3UD��A�X:OQ�	*��)��}�^7sa�(*�q�xP�2&�]��ڕ�-=��t��^���&�L).�����!�C�m��n���>�*�*�A/��,ׯ�/�/�m���C�4��[K�ͷ�As�cs}D
atl
��h�֤��Vٗ����8*���T*f�9��+�Ē@ԞZ��ʻ5�����N,؅���b�\�]j�ާ��l��A���zyK�m�U�`�ܺ���K_8@�3�T��f�xLu��A2�b��\1��e�rwk��nf��q۬�F=ζ�B�Vp�%c ��|H�.g)2�k5�J^���ٱw�]w��ؚ:�Z����)+�%:��N^^X�m��)�ho�HҦ�3x�bWϳ����@��('��,��#]��(��N>�=_Fih���U��y��R����o��������ץp.�J�
���S���T���*�x9�V�\+���$烶_�=�%�yZ6BZ*h��lxeB/^w^�v�J��<�0���T�d���E5� �.j �k:����!�p�6�}�􁣋��z��}"��_g�����ߒ �H�g5���:7'�d�2�2��a(���Tܿ	X���Q_��'q�I.�h��Զ���8����So� ;B��U_*��g����Dml@)[;��z(`����Y�����+J���Etr�N�R� �k��}\�E��Q��F)޴��']�<�@7u�+z� �Tfe�o�?aaGR���U�rX���*�D�����������ݩ�y5�o�)�;�Al���=�kf�J8��3N݉�s��R5'����Uxy���^2�q�ri8St<��4��w�㲊�?4�C���434чLD�F"����[5c$�.ǚt�q$��=R�08�nnW@�b�H�t�BDǹ�t��Ƒ1�=˽�k<���@S{��W�*9���@he_�r�*�Bf�rbNa k�<mO��F�ۆ	_0hf��M��0r7�m��z'������U?!��R�JI~F{��]���*\���n��OjJ��4���'��;\I�@O�P�g�h�+��8B?�)��Moy�����ZgW(|J�R�TG��������CA��'�|�Ale��Y�Ad3����fE���L`Hp��e������)�=�F���*^�Mf�-
�:ϻ���`�˻)�û���qj�y�?dޥ5i�(>�~<&����a�g����u˫D}uY� ��'�R� A{S��W�f���ia�$Ŏ�*o���i(9<�%�X&wl�M5y{�Vz)$�!�i�؄5%+��c�������X#��p���755������P�m�(��m���#��l�,��b>�P?� ��i=y"�� ��(�*D�
S� �R#���b�Z��;Wq,~�΍���~Ǫ���)���H�K��\/����O�T	�м���j�-	es��߭3�GJHct�.Ht����@�aa�veM�F��fͥ(�M�\�#O�xm���S�lNI`�U6�ϻ\������H,c�Z��D��d��� 2Ax�Â܈��_�m,�a��l�~�ܖ9D���.��wѫܼ�s~��/�9��&h|o����n=)`�fw�D�79��֢u��iegCBղ��Ig��{�L����x�G�%߉s�o}�2_��x����,�g�$~$w5?Ka��M�!���B�"�t��O"��E<b�=�y�G��b}�P��΍�s�/�y��r����͟<�̎?��%@�֍V�-+�k�1�b��M��?!�!`6"1Nq����ZV���M�\�sw��CSK���c-�+�)�^7K�}7��**�m�=і�����w>����xLI�� �Τ�����QkL�r�>���T�hՋVh�缏��m�� ��3���DD���@�d��5��:X��J�6�}{!{:�!G�閑[=,?>0��|qz-��t�1���C����{������t� =ylz��q��S�i��g��������*���-jSk
�����M���F�H��&�D�M����(����� e�|��eȶ]3���y�D���'���VE
�>i���jk	r[dtpu�+�]���r]���5۩���c�=!��W��w$-��eMXh	���z����
��2W��h��A�;��o�Q|�c��DY	j_���N-�|�k����o烷?���햦+�D �dv�|aF�Y&����-o*;���?�:�w�'$%��O�d���.�l@}@�_*ὔ�^Ui"��Uz���n�A6�/cښ^C�S�`4��޻�����>�9CG^bUC��J�`�P]F!�1�Қ�w�w�j�������_�{ܙ�~e]o�M�a��Ӣv6�B�/BOA�����3��3TG���R�K2�����ER��u�<LbX乗5p�n��;�yLx���~F�~֤rWYt��ɳ|��C7\�E	���!�{���l=gV�ְ�J	*�#�e1��oʃmO�$rE�
q��UZ����[oI>tW��Az��ʓ���{`8q�Gj�������wsV�,#mY��r��[Ɠٖ�U����
 9\{
@��=ꎷ��㽑� UQrO��߾��CEW	z�Lf�������������R��|�E�����34W����,���ެMZ*�����3�1�����[6#1�4ݓT��FT�AЧ��+V�'.���
n��O���w��~$x���n�զ �q�r+ً���j�4'8��5�@ ��7�:�� �ĭݞ~~rT>���8v�3��@ƿ<��Q�a7lf?�)RP���� ���#���.�o{�!\�?�k,�m3m�}}p=K<~G��9Tm�@򡿞r��đ���Aі�o���2lX(���/���4��3qq=k^�p��-�h���Y���k���B�!D��黁/٧�y�Kߤ~���cw�b������g�^�\n�sw�sVz�(����jD���X��L�N= ��Hr���|�G!��j��5�;Q!M&Kol��7{�"��N��{`I7���Pp��<���֫�by :# N���|jd~)#�'�����$n��������[�ܒ���)���5!���]�y~�y���|���E}p���� į��::�L�������g�q��.I|y��S���,��Fb�����ZY����U�����L=�l	����`炝�J�i�����}�j���P���d�y��
`xp����LS����`@����EI,�p^���]mN��N��0�V���Mu���y��x�c�c��9@H��;I�yV>����k���v�GP��{�f=�9�`�	��C�`�i,!<g��Mb+�n�ĉi��q%��JB4Y�P/q�C����� ,���!�7NZ�o����+�<�5ma����G܂���:�m�qU5}����]I�L��ݝ�Yp	Se@X[��%�W�)���O��R�`�Ź��,��{R��9�@fT�qa��v\ӏ��n"čMt�5c��p~w?��@m��3�E�2J{�pn���I*a���8|�P�-QB�E��
�J�s;��Y��%VU���&f*ީx������D��Y�����cd
�0�3�3��T%���6AU�DXRy�&��W�� �ʲ���63f�H]�8�_�)/�ݞ'n�~0�K��l4��a��g �a9%1��/�_�qI���&"�m��W�/�D�6V�&�[�D�����H���	��8i'������[?5�Ƚ5��*n+�{��i7YI���vas-���=�(M��)�PWF�Y�}<<�����鱦Z��&��\���Q����.R��1�M�v��1 ��58�J�se�#�4�X�	o��\���H[Z����8I����p�M`>;�z�pX�	{�*���uz��4Ⱦ['~k'��9\�2:���>U�Sӈ_[%���h��Tb�@���t��Y-�H(�a�������T���^c�>�&V�@�-��� 8�~uwB3dҍ���)9$�6�ګ��lRgN�'0H5*A�8.y��|/B~�C���v{ �er]E�U�q�'�̮Hҹ�g����xz�]+K�I��.��]�I)�j�׍#���8덏.=P@m�S8�����1��֝ybsV<��L<��2�~�8�6����g�3<��ھS]��'��F�&7�+�a�:��=�;�
��7
����Pf�1�K��� l�����9W�@7Q�.$�q:�vy֕(2\���"�@��5�t��k��'�?C#���e���'�|O`��w����'ҟ߇����C<��|���fo���͹��%fb.;��_`T+�J��I��� 2������Yy?���Wߖ�N���l�C�=����#h>���Du���P���'%9�wx?�);�/�Uێf���xq�U�}
?�UT�U�^�\�����ԄgP�f�YiR} f�d����vlP3b&;�?��CU�=_�g<�YE2�nJ�O��;��NoD�$#�V� \Y�S��`�����ȓ��������Z�s�';���6�����R13���!_����
f��MOh���W��Z��Zp��.럠�g{P<sX�b��=�CY�/r�ib����O<�E���qi��4��R�P*��y]�I;o��*��z��vC����f�H�հ<I4k*���h{���1ﰩ�pu���s�c�2[S��������W|���/Q�-��nAK)�}� ���o�7JߖWƒ�,�h����[�����J6	1�-d���d˃b��6�ի	��@�u?��ޞ4�ِ(F&?ꕽ��'"�=3�[m�0�.���ѕ�t����!�ȫ1S�
�s]����i�7I��@`ߓ�=��
�αZ��p*ƦZi�ܿ�Z�I�j��H�lۊ8S�#z[ݭ��K}U�چ��̽θ�$�|�؉X!he�F��K�(4�ug��'(a��C����P��N��TuǏ��A���#�Ų8�b�M�'䰮��a�0�� ���؈�ޕ�oX�ZI�������)����W�i&o��On��C�-e�CpA��C�����T�ʪ���z�6Vk���7
���Ϫ��g��� �@��z�;h4�i?�E�ns���QT��ett�Io���p>��r'�9�6uo8xC�~9I�G���Y�\z3�9���++�&�L��AaBX��zP\���O���̍v�����z�f-ofn�:L��uÿ�)��r���ވҏF��* ��uP"��1���Ņ�ٯ������t���ͪ`_E)��3��eq����7YG1����<�q��ҥ����:�Aq�Y���ہSt1vN�.�(��j@��Ͻ��>��h<G�K��t��*\�CZ��0c-ϣa0GS�Cϱ�x��ѷe�Er��Ey{Ax�M��dˤ؜@�唨��|�!6/�[�$�9+�����=R?i���U�Cc�q���c���}���IC�L�1&˛�y���ޖ �z��{}Wd��J���+�w~��W�;U��-!k9���9i��N �Vӄ���M����E�C���[��ݗ����%�Dh�����ɓs�̖����^o�4�
��I�Uz�Ƒ���M��T̑��u}́{�sY^�=>h�27�L�+�f2��Ĩ{A�Դ /��P��F�s��מ �k��b~)׾�ϩ>�)!��?�J��=�[�'��ƙ>��c�S��I^��P�WS�iG�"�Ec�'���V5$�C�#��dJMӖ�^�!�5Ȉ�{f��q���0(^B���\G)�$c�]f�7)�|4\�Ǵ�xV�I�5Nk�4?O�E�Bv�Q`�k�N��h��O��GonO:�S��w��'6�!HAl��f<v=�V�n�IOBbET��]U6xxͿK���0�39�A~��N@�dz�����^s)�珸�x��~�8X[b�`E��;s��J8L�I�o���;Ov;�w&�A�+?��ߓ��N�m�8�(~9�g�����qqA��X�vb��
w~������=�jr�^��� ��4ݯQ�N� - 8�$���*,�6�O:��d�&�c\F�G׏�U�U�F^ʵ�-C�e�_^H�V��|�c\Va@"���{?0��%�xQ]��é�=7��>X`\sv�ߴQ*�5���S|o�]�RDŰQ���1�3w?41����Y_�Ǒ-:Lj/��tU���Yȸ��A�E��7�Ɉ�fA��<���PJ��fz�ge^2a�&�6/p�w5�P���l�y�ҫ;�*�nIR0�Ӊfmv�B����X?'��_�&� ֘`�.-�S�#��&����j@���ź��7��]NxWث�,��9ѷ
l���&wM�&e��Ȑ{��X�_U̗������A��RJ��A�a*��%u!���Y{m����"c�g'o�RӾ;���`Z]^��u9kV{�Ogq�r���[E.���2��z+��WUHzR��x�I�z��#�r��J��G�u#%"go���Ȩ&��+���Vt��V@j�/;�$�Ԑ�3�B�5��+��m��O�Ƨ�Ch��؝ˢ���Cb�	�{���
,1�>��b��i0Tw��?2�<娻@K���e��-[���u{gx�r�CaUf�m�iZ�hF��3�視"�6q�na�Z���j7���p��W�!O	p�@N�L�f\�.��qxi�Rh3�]Kұ`��j����z	3^�s��XFV>"���@�.f�NJ�c�	��ާ҆�t�p�X}��}ٗ�-&�W��Z�yi�E�~�ػz���u�K�T#�$,������� ��7	��S�
=v5�BY��S������+���	2	��̐��j�D��1�9���Av����F\��Cs��i$֎�]p�4�����!Չ��N�к��Pj�c��jL_�6�d��y�X��&oX�9(�!V�ے�*8�;����]�`�]cԨ
�P!��*��12��6jZ4�e�y�d����+�O!�M��=��>3Ok����X!��{ �{ק[e�L�^~��8ND.�%�[��ܯ�y�&��`1�#����O�Wzd�����#K{�[ �4h{W�P�{�F����&�^ ��O�ͪX �cs=���7S?z�"lOvY�L"��!+Sˋ�}�����.�
�~}ut�����n���w,��x�0r�Ͷ8��H�3�Wç�s�b^L����e��:�XX�.��h�'��s,�ki������ܒ�Nm� ��C����f�xӨ��v�(j�m���Z�$\	�PIx��Z�8A�g����g?�.�"Ͼd���HA܏�h��c�K�U̚�p�`>���Ա)0�V�� .�/��EL��s�V��	�l�����J�D��/	x�����HCBI��� �W�\F�1�AK�t0n¯!B㡇��P�ڃ��
�����J����2�3������ÛO����$`���\�_��w��t�-�f�d#"L0!�?�\��h$N����7__'�h6�K�}�{�si�9�������L�9�%s'<�������P�𛴴Y��+��Ì���z|	O�QP��>�b`�e��
�!,Oy�"�m�-��Ҿ���|�.8 ��Q��<�p ���t���/������/��63�>�H�yʯ�ٍ��KO�z�˙W4���sY|����
F�i]dw�m�s�{Qn��$����"t����/�L��-����8��e��}`�h h72�8�/:~�_k�ֽ�U�����S@����m!�z���q?:��|��B��'����$e��W�w3�;�	��Y|�ɰ��H{��G�S��d�	 ��T#����������r�e���x�I6F��c�tt4����7a�,g$RJ�)���#xE� UyRo�f���H�3$�r:/X^	�?�5�qx��I};>u;�m�@gǦ�yj���e�0��ϫ�}Q��^�������q�I`���J�@�|��㣫ؔO�������`�];h`	1��q��up�[`\|'$��3�������KUD���'�r���<k��D�n;�-�����eE��r���G)!8���B�9��{H
� ��EQ�m�pJqG/��l��x���
ϱ1��8v��~�m����~j�"��I���n�B�E���q��Sw��u��^��h�`�g.�+b���*T�Q�yMN��x@\z�V�"k�M�3�g"[�b��D�lH��Y���u�~M�8h�S ��o��,c��U�Xz!�=׻8�B����Z����n?���kIt#
���Z��n�-�j�� ��w�xa
gi�%o<���ϣ�����<�w7�#ͱ]�:_�1Fى��>��x��ͅ�?�뉆���d�B�*g�։���P��t�S�X*V�c(<�Ԍ��(��5&�`�޽v�ם�W�a-���>����~<��%�$��1Q�1v�S������b��ŵCn�D�"	���l���L�� �[��%A����p�¶#û�v)-��>3�P{��|�]	N���,� gŦ�
(��1�8_/�T����g������F~�#��C"1X:Y\�{Yd�US�¼�*��U�����xΨ�e��I�Ѷ����`Sc�{{�'ė�~rr6���¤��5�2��B	2o�Z�.7únس�xzM�A��0LN��Ky����)����׫��?�pg�ʶ�|���~�>�@���}��k\�=���;��'4ӽ�j�Q� �.�Y�gL|M�ԲX�N�!���� ��[�\���U��א)�����/s5��?�-���G�s
1I�V�i����ì����D0��e�܍�Bd����CV�G�|jH,���a)�d�.8%~�{y���C�ڹ�AK��s��5~�eKYX�p��me�n]BM�X�ǚ@ư���\���"x�������N X�AuX8t6�lp�s��c{�t�����dg��F0��5M�-V,齨��y (t��~��EI�1
��Ʃ>��`�g�݈�(��8��D�*�e�?�(&;�Tp�H	8���R�(� .-�H�<[
�P��M����6�xh�X��������1f�v9p	m/B�Q�����	+ ]�}67���=�KB9��Wa���l ��������a��<z9@H?������ �K���޻�3��3�>�<�N��T+��F f�X�*ݘ��Z O�Z7>��'����jl���T��ND�*PS�jX��ۆ�Э���A4��M��;�M��Ћ!�nq��lS����*����%_��� ��π��F���mvU:��QU����ý=J8�`O���6���;
��^ʏ%-h���v�������:���c]M�s��[7f>� �c��S��F����y�6� �\�����uT��ݩ�r�yfiñ���F0wK���Rڝ� (MrO��NW�*{��w]��ҥ��7$�����͹F#Kg#�����~���C�T ��!G����(ɑhN8������aT:H��*O\=K�ѱ��7/��'���p�5�
߭�F�rG'�&�]0l�t������ɶQ50���L7�s;��ήIz��iK}r�)6V�n��+n�_���v{�[�����߶��Zq�P=���jYf�D�x0t�j�s��ř.�S���s#/h�$5E�9�h���K����B�z�0F_��{�)����V�~�V~48!����DF�մ�����d'=2_;�K���������q��s�S��p��*T�Jr���W�I�)���p�\=��CL�<[3�A�		x�h��}�tb|:-Ł�~�Fъ�k9/�eD��I3����4H�#Ǐ-U0Z�g7��\�S�3����ǐ�|�	j�94���r�����0�u�U\�$]��h�(�*e�;d��<��G�]|/ᇸ�x�&���Z-�𮀐%1|r2 }�����g�-�T4�b��Ƕ�ۍ$�@�Vj�[[Y�r�4{1���j�n�-#�#�dN�u�d��u��� ���!��\'���PP�=�S�͢.��Y��-4P�KN�z
�tR��T��K������p�V.�{q�,�<v�®H�{�Z�����#�Ml��b�i2�f���$��d	��%�m!�az�U5>����)��N���r}kv�i�Jb������ô�{ v�]�R��,'эZ�*Thv.�z+p>i=ڛ���G�����S�_2�0#�;����;�<ҥ���O�'Q�5�D��I��q�>ާ/����O�n������m���B/D�T?a��>����3�M�t�K@�L��)��?�Y�(��`R�L�|~��S��
��1~=aEG&�n�!@{�~6lI�Aλ�����1�iu�����a�+���~|���	}��o��T���ݫ�KW�;`�z@5G�]p� V .�yk���O��F���3��D��\�����k��&V�:o;epq܈ʞ3��A�C/"[x�@�|Q���X]�M����Fߜ��[�h�H��&z�Д�l��?�� E����v?x
T�V_eclc��B)�_l�߼�:aW�Q���)�*z?�:�r"��g�E)�T���:Fώ��
F�N���ׇa��ߑ�컻�ɈK�DX��p�AJfN��ڰG��(Z�A(��Fp��9b��e����}1��3��?��zvd����_`���f���b�hdniЃv�KùԆ���'#�o�����a�=��؀	%s�x�a�G&�os�X��$k�'�Pϯ�uc����ֳ6Oi��J��]��T7��O1�^����w�LA!5�,���X]�Hn��Ñ�S's�{�t��5���5��p������F����k &�����K�P�XMsR �z�$���v�Ć�ܻ�s�8˙L1 ���@�9\O��|�[$ �ÿp���G�f|��G���M.��ܐp�ѹ'���3�ŕ�XSyCqޚB�q�m�P����l�+�8#T�Z��]�P�"���6��g����](���[ZLKkP���oL9m���¡y���p�x�ү�(�X�x��Y)�3,T�����I��W3�G�*����X�b��\��ݨ@ΧuW7�!�*"b�gq�S������=��"��w,?�7�&�ȍ<����_�w'�5�{�U����--���ݣ!�듘�;�.��X>:.�2��'����L�LK���������cޱ��F�Y4"���~�K�I\LhT�S�ë��>���΄G���	������U/Y5N�s@y��>�/�A)�`b����%��S
i�\A/kSR����L��R�����"n�����/L�����OS(�It�)}o5���fzF�D��c��a͜��>�:�a����@hSB))U�=e�+'���Q蚩{{����y*���){51�Z�:�,yl��|-/ʦ�y�τ�B�O}��l�J�Ju�x ��A�S�ɋQ��n�l�f�*�
�Ne�>[��*���� ^�ݚ��'�g`��s}�"i�lC&Ӗ�t�W.jܺ�6
xv(h6���I��$�\L�������,�)�HB����E����gVÙ�tp�Q��>@�j�����/��^m>� _����Dp��! �ӞC�����ܱH'�����Y|�"H?!���w��_��m��w]�˶�i�Br��G�|QM>;��R�6.���}���w@�b��~���\�b�g�䤪/[~`e
��C*Cኒiv��(ʄ�m֏��PԽL�����R �x��7	��>1�@���d
>�m%*{����j�5%GugKf$�s��)����_r�8�#�[�%���Q<_Y�7<"\umS���-=YsfO�zE��T�po!�9�8�PN�2��A���C4˞� &z��~`��6y����V��{�,�䩕��9���$[d�`���*uE���������N�&�>��T�`e�4*�a�6M�>���h�Ϭ��0Z,���N��W��!�,P�����
jr�~_�F��[�6u���z��&�>@�S�,�U��M���'+�|�F��45kA�HbA�<+�@D��c������*�oBp Ͻ8�{Ὲ�&��g�:Y{�'��r��u>8�������^�:��pĮ�L��Z8�9M.���ΎgT����hD���6t+�l��ʥ�f7&>\5,���s�����
�̹��Ô9e���O�����,v�D_*h'7;f *�3[<�ݙAckc�s#5,$�k5�pv57X|vh�n�����(��{�,J����F5�D��S�����	��%9 vm�+�i-*7X�Y\E�bni�3yNc�ܶ��/")X
�_����8+^=��Y�X�̠��4�m
��m0��k��] �6p��K ��c(c���ՈV��҇k�Ѕ�����2�>�2�`���oOK�bcE�-�^c�/i2a�۠NT*�O��шP�-i����c	�ٯqYO���R����O'o2�?�W�v2M�& �*�
�oT��	��kg��C1�o��g�:�CͦRVa���M����*R��x���x�v]�U-�����:>���i�N+��Ke{W��m��~����!]YX9s���d��E|ڹ�z
Uȶ�R��u�>��x�b�/�
懎}2�"r�¤Rݛx�����oEָO
x�e����ƾ�y���"�Kl�w9��C�͈�E0g2�� Ѡ�(U��a�TdH��>�bE9��喴��T��Poo;��a6����[��Q���ؘ(J;��A&��f�GQE�O��%��
����-֐9Է$V�H�釠�.,�z��T�5�
%)?����(,9ѱGiVQsky�f8����#b>��=AsY���,�n��S���n�d��;����%״5�shi��	���F��t�ϝy�ֺ�����w=�&�H�f�_�3��?h�L�u	\*ÚrP������h]�Pի��s�;���G��gk�<D�xS��t���mC�M�֕��;��>�R��BؐLְ�|�w��1��V��;Vz�sѷu���= �w�LR_V�M�T�k��;�i.�?��K��e���~���7������L4��i���Ԇ�p��A�E`�R��GK�Q3��e�D<�t�|L��Y��)�4��k#�9�Y,����������^�9st���,�0vZY�ģTnX~�J�Zv��<���aJ��e�3R���Z�����#1�R�a�I۞Y0�Oz10�/��yK��V����fꄴ[5��<U���+��J�u:"�a[h{��|(�Èkg�����Em�8o%���XŌd�&V|���8�O�k�4��V!O��Egw��� ��������x�%-vy"V0'��q���Xl�T�ћ����M։�� �!Ua'Q�u�����kT>�Fvo���
7�4������M2��*$IAFfmY����j/Y����)E��Jf���.���M�P큠�����`�h>l�_+ϛ$���ٕM��6��GRSӧ4���O/$��']�z���Y�%FX�"ˤi�@��NwIs�S�8��\��A���Gb��� �w�_d�˯�:�Ň��Gu�3��iHN�#oH�E��/�B&@D>4M�RA�֙��B�uzKt�	M���Z;���rì����*AɊ��r&�.��
��.Z�,�3{Ø��,$��.	�����h��Pv%}�E$�4ʵ%N��e�.��XF}�O@[TbhSrD�(����*Q��+����{��'"��j`!D�D�};�`28�̏��J�W{��%�z�n�^s�
��@n��X̰�?�)��vi`�Z�B�+�e����k��i�5G$y�:�r&b��W�=�?	�^r|�����͇�������ꙵ���3 :�9gcYm�R�/q?�Lm�P�9K0�)���lla��!t|�w�����!�΁������j�a/g���WP[���b4hu���KU�z������.��`*��'�K�!�`I�(B\���H0ۄ _m���Qdw�����Q��x��e �X��D�!fP���m����Z-��Y�|�wO�I�����[T�6�'�^J�,��Y�7���<Zӛ�~�z����:?���ڿ��n�J0�03v��\��Ɗ���U^�+n�@G����)�_l�Fu��w��@s��pw���
|���P�.�Vp��$]$*�:ܕ�pb)�1��7Ա����d�ag�[�Ke��f�o��hY�+5�W=�s�6�׼�ok�:�:��@��e`F,�y�^���L�'Vu(>+qj�y��H7�8��fϮT�M�o�t�_e�:-�e���8D�
ƝH��6;��_Wق�NV����=��lw��|�����N�0�[&�c���"����#�
h���oϏjp�
�^֙�S~�,����Po8��IQ�(���²Jc�r�dvY��l��Z�����m?���q��I~6�t��i���[S���GwzSlMp��نr>��g��D�qD{�l�5�5�#z��j�	K3���(LRp�KT����t�M�q�����'�I'�r;)����N��Ȑ ���'#-�A�o� =�P�):��Rm;�.d���`8v�*���/%M���5��#A�C��*rіvwF��K8��_����Bv�����A䒃)yp�c�J�	��N�m�Ӟ��r���N�����Ei��>O,�c�3F�T����#mM����p07� ��������L�g� "\�}�R �.�2�Q�%d�r1��n_��r�.�0 s�7�3j z���HsM�#pZk��!si������=�Qu:���6O�ܡ���܂u���ɬX8��,�|"���?���	���<�G�z��h�)��5�3������[�,	v��؃�d���q�l���F��؟�?h<j(�H'�TR�d�}�y^�G`hBem~)����="����(�E�)����:2��A%����h�!���ZZ�(	��Ջ���>��`)jPˁ�����b���/������2�4�g�v,5��y�a_����7����:B�jA��d§��f�Lp	��X,�x��u9���M��:�~�n2&� �T�מ�V:�|���1jJ�0TߚAn^�Y��i�,+g�=��EZ���Z~<� �c��9�fN0ΐ�U;�%�\,�p��FzY,�P~�AZ�����Zrvt~��+W@�{��~bJ3K�o�g��@�?��:�.�E�y�0��Um�0�U�кu�EKH��&n��Q{-l7�1�4U5��@%QG��/�O���e<�Ӫ��:䇁QP+�$�=.��;üx�bK�@�t�YZ��6t�{�K��4��3�C���k�Ѻ�7Ux����9���[jP����>���h�p5.9ϣtz�;Б����D6�l��W��Z�%���]�1����ȅ l:��}�!�kfO�u��q7��LͧJ��~�P�Jsrq��NOC�$�1��k��\��Q�U�c�?ֆm��גKꗉJZQ����k}����Fy���t�}�l���7�������0'�Ř
KkB��:]�Q%��-���Q	|f}��xJ��g��<6d#._��AEq�Lx��}Ei~Q`�a�b�@��"B`�A�� �Q�~p��p�Xu7�ۇɶ�͓��Ki/O#��S����I�Ȍ_����&Ǎ�˝z��D��j��"Š�xd[xJ�勷ˡ�#��������m?x�o���]�.�U�3�_]z���,˔0ݗ<��ݓ(�=Z�9-�O��^�h)���`J��xu���VC�So�B�p�k�l� ɒ
���*M��3�@�l
Q�����S�40� �OQS����������V� _V�S��V��+SU�
��whp���ܜ��<��(V4�
^0&\�x�%���xz=���C#nC�y(|�B�V��b��š��C�)�l;��b�> �lU�;ޞ�V4���.�������0��HV׭�D���b�\��Χ)7^���&�[�H�\M K��a`��c���^�)�խ$�8�;����r3L�7e�b[�.��|k�7�v�\d��A���S7"f�_�v
5�iP!��ѱ!�s�]���q��w�Ŷ�����J������7I&�e�I�M�� ��k����Rl>t���{*��HZ��L���U�v�|{G����0�Y�&��[h�l���%�Y�P�>
�{��cZ�}����f�:3�-�tI�F7/�^��%~�W.�r��g1���K7�e�扬�^yS�jx�Ơ��������Kv�X1��b����x�v���
���ye�oq��s�5R���b�y��/fb��N�c��)����l�����-o�:��(6Ҏp���B�&���5��ɟ�<���6=��P��[У</g$.]�s0�ͤu8�J^�~�`.3� i5�u���`�uS���kB%����`�@u��#��y�b�ލ���Hl{����@��YSU�y��2�A�R����cPx�y�x*]tr�#b��N�V�4�Y^N�nM���&�Sy�+�?-�訰H�[UC+�b\���]�u�����YKn18� ����ie��K{��M�}���B8��\P�?䵪g�����{�iY��zp���'�0����!_�Mk�>�G�X��_���Z�g@�
HȞxw8��X8t����︝�(��J��}�W�m�Md4GlԞ͊f��f���c&Y��܊��H�2��o�������յkB�����^�\?�ش2�/\d�*R�Ґ4���3�����Ry/�(�C���i�`;�0�[��5�޺���t��_�~3Bi�5t{N�Ri��>�-P�a���d
�A���JW3��ޡ\�`� ��3����w�;9]�a5ж���a�^gJ�r�j�8o c�9�!ipǰ�p=A�A{G�w���?�dF�0o�#�]���=c2���7�x�u�=7E[7���0�#"xڷzrĕ�4���әq��f>��W�3���5X,XS� �Aio)�u��4�y��ѓ��/�ђk�|p�����2 <�g�[�n�C])r��$��|�����}�8���_���t��V/w!�[���kiȖڤ�'/t;��@w{,@��_����v���b�������){���c�����b�g�����ǃ�\���`�3�I&��%� +�4���ylZ\k�t}��U/�)�:V�'I�>�{ ��ȭ'�q�������~#���O)8����ӋJ�T���'|w;F�"B!�0)��`�<&�&m[7/�v��}U㑕G?�X0		�G�pỲe'
�a�H.L�Ԛ�$G�۪�檄�DU�/����4"}I�W=*���8fz��!_�����I3���zW�
jw;Ʈ�q�fźV��i��?5��'X�I���{�y����4�ha��G��@8QiE?hIK�ov�ˈ�<-M�L��"�R���[�����?�����ݍh>�ZB#v'�"ٰ��ߤ�I�e�7 �C����[�� c��9���^P5P��e:�ņ�+k���є�~Sه78
 ��X)mrӮǓc`#��t�[Z&���QX��|����ۧ��������'
d�0�F����g�u�Q�j;ŭ��2&a�a'޻���Tucs������QYy�k�R��0Q�w6�%<��u��&��[��z�L`ٯ�-7��� �ݼ_�?O�&�Uz�s�~O���u����B��{%�4�U��O*�W��E]	R�L��~���,�p�z��U9P4�6QNh��)6W��gw]�=�OB�+4n�?�&N���� �^b�h�zQ��r���u<7���{��r��?Q��� WL�zfȔFv�8�,��:� '�Y5"�(���ۢz.��1��GU�3&�֝��1i{`�R�}�6� .�G7�C����jf7��]�S�{�;[��^D���}4^\���#��+1�w-{�0�^�@�jP���i�^�Of�������!H��ޛ�=`��X���/(.l,���;�g�5'x��-(�%V�wFS��HU�^����,^�<�.A]4�QC��4�
U?�P�><.)��`�B*���$�n�^���2�p�&��j[��V�<c�
A�X�PA��� ~���_�������	�C���Hp#4���'В�ՃD\�l�U��S���n�5��1�J芃Ke��T�(7�G����}��Z��<8νQ�	�����Ι�I��FZ��?�`��5'Ge����%�Z�Rsg<p��?p�iaۃ�������Nl��2*�c7�s��UNI��٭�������f���uW���59��6���U�Qϭ�sS���ɮ��MM��|-��4ޫ�*�k�=��I��J�٩_�[4��f*-,��I0��x�[�&�V�ѷ�_\�$fC�Lw�P��w.���V�	�|����މ�3Qыa�U�rʣ�G�����[T�7���O?:����$.1��E��
<) �}Ԡ�31$ e�(��Xy�ʍ�Te8Ւ�Q]޴���G�.�l�kO� }��|3��� N�[���	�S�<���Ċ_��Js��;ތ���|m���T.���-ؐU#IX�|g�D�C	����Wő.n��-K{I��j�ēϽ0}�+}�_��.
j@^m徘!�.� Jժ��ӱz�b��GM��>�u�v?��!BW�L=Gw�lڍn�Ft�c%(�c���|13y����г�fשu���"Ë^]�	�kP
�BWs1w[?3�Q��� ��Q3�@l���d-^7��y�l�	ٺc��J\�S�/�$�]p���~`��o +����3�<��&i
���i��������ז��
y�,���gm8I�i�qx��мB�Aa@m�Z��l޷��=��Lsz� �k[�Kt��^>$�uI�G@z��"`���J�e#8��d���b���� ���>/��g��RhĂ腌�5��+.��Y�rJ9�$]�t�淫�l�kZ{����p0���ْE�����S>_�nZ�0�9������c���.A��_V�;f�"�XyxIGx]��J����KQ,�`˨u����Lf{�y��G$��B��9�*�鏎oBd�o6&���N~����r��B��s����Wa�M�z���<��~4��a��d��5*��n3{��^V�����e���31��=��%�PĕVwp�c8� mȌ��U����G �a@��*�!�Ρ���2��V�I�����=�܌)�����?	�H�l�y�?��a�t��S��/`�tx��L��T��<�H�x��.%��Vf:s3����zٺW���ԳQ����¿虡��C;�m�ʖa�X虖���ab�<�m�m]�g�\*�Ej�J�I�ZS�{ȓ�)v�^���P.��1��6��-.��$ՠ��?ll�ه@R�=k,	Q~�q?va��R�|&�T�,���\�q<�U��9�rr+�h�*J5'�.��l}qM����z+�Q<k
J@5`hظr4ڴqVG^�������u�fxD�X�N�eE��3U�,��J4Jt����t��A�����؞TK �
�)�KpR���!��W�%⡓o�E�u9��3����1���&K� 	Ej�ߪ��a��W��-G	��}�H����4��3���f��7D	J���������`ҁڝ�V+��bO�t�j�r��}	]��&�2_S��ʕ���6��sc��h�]n�7Et����@�t>& [�0���6�a:@2����8j%�J>5j�vN����� w���Y�r�����w:tE��Ծa�ȯ}�P�^�r3�&��	&H���x8sv9�h��ɫ�5�K.U�ۆ�.v�_W��cQ�"�>7X~��f'ㆬT�=����S�̵�nV������
�l��*!�!}ĭb#�:T�^b�&�2�ҵA`�E�F�m��t�k!����?�mp�^�������m��ѯJ7��~e�)���T}��K�<��Vf$9�FJ�:�4D_q�w�2����ܝt�I~��j�,��#(�,�l<Q�������1��N-ˣl1�Efs�`Ӡ���7)t�� �����������X��_�}�۶<u'���Q+u��z7��#��X�y���W�>3�Q�)��WZF���n����u$pf���|y�NN�ZPm��ǽ��g"h-�W�lqQ����` o�}���'�1���?�)���� ��>ɤ)`z��� ��(0��~��N��	�%��1d�}��3q���gP,9<�k��={�I�Kv��1C*a��B~��b\u|�rM�/G�u}Õ����2i�C)�I�s1GTļ��-ЍUm�,�� M#M�����
���(�8�s���"�^��@t_��e���YW���vL��UQ�����]�Ur�|,�pv]Գ����,����ђ��=��Sشᷠk'�kЁxVZ�>G4�L�#Q��U
6���R�2,b�Jl��/3�� ��O�F�YK	�s���(𝌵��5����̟�r�9���_�N�R�����'O��h;�]�<�
�Ra+K�)��.�]/k[ŧ�D�]w�F?��d*���RWEx���Ԏ2�m�[��|5��!�g�V�3�l:���Uژ.~��8�0�W�!@2B1���]ʥ��F����R�ejeCw�Lh0���e����V �\xx�`c�X�1��3���2�z�:��ߎ3Ct���=�A�5��	�A����-�C�s*����:B,�9�8�%$w\Re�k��ߛM{q_8[�NL/���`A�('P1}2�͑�s ��ܚFf0�tOfr��_�g��Y�9�@�ezL���I.5��h^U:ȍ�a�^���E?�>GӋ����:	h�
G���tC�<�j��tH�C��c���Z���4�=U��XZ�
�H��5���V1i*�9���q�-����2ՙ�浱�;�����-Sރ=Q���%)�^�|��Z�\���ou�8���:� �k����r���k��ݾݟCA�C.D����O�/T�t�����x?������pZm)m �8��秒�8��ܥ���Mj!�	��š�����vy>�Ŵ;�>��S�b��Ƅ�� �P�$�E@ �����Y]�1)W��h<{������Y�֢�Jk�isj��fۤ��ktv����l���P�0���GR?4���8YV����n������I���r9�E:�*j�=�` $�]?��5��C��i
��#5r��M)�c����%����Z��aZ[���T*]q����ڳTF4Krҝ�
�.�v��w�γ�^����$���Q���6��,�z���^��q�hɹ��X��,�k�\�iU�%� <�K���`����v��Y����/H㘗�.�����V�Wv�˰)Vįz	s{蝹B�]-G���F�ܳ��7>_��oA O��*4%�����2��^{9�.A���^��Yo�&�n��c�g�6h/�"�����*K�Rҭ(���["�����y�]�?��a\����	ԭ��>��:�]���
;]�x�l^���m-�T���-�~^�ԬZ�Ƙ��b���P�F����Z�XM�Z^�H>���37M��R8��s�M��7Q���
��\B��Ϊ;�%�!o��ٹ.ＸH,3�o�.ط��½u��+���>���ᱵUQ%��t�w�֥��ÔO�G�1&au�[L`�O U�:iM�r����L�<�� V�Gr�u%�?�]�:�-���	�sj�,�J��j���(�e����몘��Q��G�D�j�a���F(���I"�M���������}֗��BE��?�� f�&��sO"��-k�>�Ц"�3��Rj�Л)AF�[�������Y<������˷�a����OP�$���5�p_�ʑz���/�E�c�ϔ��w�x��������nP�4�s��y���{'�'�^�� ����Ӽ����.�>x�k��3��@�^"�>i]��R�"yNQ�x�&c������$jl��g�[���"�,q�p�홝h�I�Φ4@bc�.{ZON�����`J�!B��P%Kc�{��X2@��Ɩ��#���v9Y0���<��D۱���7ݨ����4U��-`�f&U�]�ظ(�Q�p���ƌ��Ui�����H��ۼ�0-�] �j3�nvm�A����r�v3���_ZSSw��X��UM2�+�⻬Ꞁ��@{C���)|�W(ho���K��Ls��;�[?YءH�z���SPAz��aX�8)���J��ڼ�8j�B���~���%�*�]�2���%_�;.�O�����J�Ry*
���ѵ�*u?�j=�$x`s��؊$�n�`�-'V3�8E�!(�s,�Wj暕ߝ��&~�!�["���~����*,b�������8��p�6�o��9U�� �wlQ��Ϊ�Z�)�5���l� �j6���Esig��|oTG���4W~�'�������'��؃%!O�~6����zh=������B��]%�&'e�%i���h���(�;��غu8�0��.����?綖P���O���b:��[s�N-S�HPw��+1�H�����9vI#��K��yɔ��<� �5����L*o��y��X<)�^��^��ϙ�\��x-c��:i��4����3�͟61�Bх��!�����z1��>����md�?�_4j��$��4CsWk�P�r	�dq;��ޟ}��f�*!�#��
��Է'�[X��DcY�T%���9D���.yMJ^�e|���BC�_/�/c��/ZԨ��@��+t[�C�ղ~��k�o�^=��	sh�&W��k�� A�B�5;=lʔ�!�9���u�f��s(OS�n���ZԔ�D�SB89"��M�`v,c�Mb�J���"+Cz@���N��ƫ��ho5O�s_�^�� \:g][D��Y�p�����K��G�c�l�P̓�mc�3�V״���zD#6�G�E�+�VhL��3�� �[#�O.��?�9'�o��A�l�@��u�Zt�*�hC[�:8�:8ȑ��Z-ۜ�YG�u<"��!�}�3�3[a��F3�`�'*x��'_6.�@|�jH�����6'Et����A���H(������s�H������<n9�լ�k��� �A�_�y�ʩ��A���y������R���Z��F��r���W�����3���Ȧ���O�-86��0� y�Ɏ��Gk���i�bE�?���Ha��û�?�V��T��7��G�̾����n˟5qVz�{VC���.���6�vJ%���aP8R��W��JKXne���"��9hH�5&)��)0�	E䂮x�6ޟ�c�����bܯui��}*,�i��Ԛ�|�{��tkŚ�!w��ڠ�t��'N�n�N��?�{A��]v@���Z+X�\�(﵀tE��;3���N�֣��*'|u�j�.i��!����
.�C���H��O���p���9�	���!��D+Yoܤv��U���6Lp�)��̓�p�Q��uR1.D�$�dI����6�mCUX�P.���9O���{T�䊹���O�*oeƺ�yI�����>���A[%����mw���L�Bs�򓎢�W�m���J�����-�o8ä���d/*#�����K��X��;���Fmd��A��7�NEN"��r����2����6�GƚS<it�b���9�CX��֊a/��g�|�4�N���3�/�	�w���o��������"��2�2aV�d���P@�Xb�^ ^���������?��V��� �gE޽R�c	�T%=a�*G"dDJ�����?&T垣k+HW�A��/��m��`ݗ���B!sm��r�툳B��K,�L��]=��?v�i���۝��:d;'��%���W�[W|K�kgȑ3X�^1�<�rI�ZM��MU����V��n��Ҹ�9� 1�r��ﲦ�[�dtz�3F�y���B�U+z�ؘ2���.��Ø2���e˺�71���pϖ.T�g��k�{,�HӖ��j�3���ʪ���%.�lT_�)����>�T-:yDƞԎ�򌽃�������= "�X�O6��^MݓsT�Q�	9�ZC[S��G��������w����W�:n�8�1nO��%�/&�	���<�s��u��򆙛g��t��'N��{|� M|vY��0��~��)qƞz���g�jMz	�]ݣo�髅%�%����j3k��7�{ӧp�D���Ft���� ܅��R���0~��q��Ʒ;0����i���v��2�F<%	��F���!�BYK~�Zq3M���T<���g�,:�*�������PV%k�c	�V���s��'�(ΧL8�9����$��bc����sѫ����7ʺ��+��ܼ�bՉ(	��u�۲N6AW8��傖4�'�D��M��ɯ��0�w�k಩!���\�3�.�S}�O��t�<�7d�7����$�cH�"PPc����-e{py9�U"M6\I��^�e���X�ˈ�^l�u����\T�Z��8�R�m�:.Gk]�7��G;�{2ͦy��~se�+������jkƖM�����څ^x�����B��=�0
}���i��[�)�x�����:eU˸T6~5��3�'��_��\I�g��n.�s���Xl�	m��4H_s{���d�U�r7�چة��n+�i���C,��1�4���3|�*s_A��w���3.��)ï��f�CV��ބHq��~R,|*��/RH�98��Fͬʬ���r���s�U��,m$��Q��n!�1���E���LE�I�����.R�����"҇U��4=����n�n$��<��EV�(th�i8� �}���X���M �aj�23:
L}D8�=8��!�	��A�'�8�"��)(ۅc*��z��Z� o��Fv:Tq�V&fPM�ƃ��f8O�z��B��t6|�RWy�N�{{��]���]6b�����d�/%\<���#����"���"e߇����LA	%%��۔xkz�H�]c+n��~4��\Xo=�]{"���(eY��Mpzt7TM�?y�4 C��˄?�OV�y0Z�H{�wL����h�-[($���{���x�_��2��P>���)�U����p�%����<�!�^��(wqH��BN%�������ƒ<���!=VFt�7j��C�`�c0��O��h Er��8��'�B�w�Ƚ��������vf�y��MQ�Sr�ڏJ����/ش�����/J_� '�n��]׺a���2��Y�;!v�t�S��\v��rA0�*��eamk7�q���{�b\}���j�qʶ�G���`�Љ���(�4����\jjU/��p�ڟ�ܭ�Ȟ0K��=���
��i`����#-��e�h��Yx�����e_mRr�7x�����ñK�������m���o�w�fM��C]�W>����	+:s޲��<�Ӓo�^�x��S�'���sx}�/ ��bRw�7~�e�Ѕf�q�¸�Ǡ�0�~m(dd�<��`��w���!�p�����3��p���K��VGor=>�ψ@N%�i>MAX��˫�d"޾3,��_��/����Q&ԡ���[����K����ep`��(�?��dW���ߝߨ�Lx����Ζz�P��C������=����a�}򄇯~���C�d�����k��ꖖ&����$��T&�,�mN6�rIT3�7�N
��+��RP�\��L���q	�(�>R���F\�����6�Eg���H���iTfg�ѐ��B�ӵ�iL��Ê�u��W����x?'��t�+�kk�Q9�I���1�F#��*���n��-T�J�����1�0MX~�ӆ2��] 5��ۥț<k�*�Gȭ�J����veU��ޥYNI�(�n��z���>�fo�&���a,�H�^W�K|���)�i�\�h���:LB��:�e��������n9���	p�Q!�.=*G/ݴ��|�klC�Utm��6�U�.�<��H&y�R�I488o����	���8�Ʌￇ��m�|�~tL��6�뉹{�� ��jւ,.��vv���m���� ��hƟzͲL���oC;�ز&&�o!�)^ݠ�9L1��!�e�3�Ll�*e�T���"���Lu$hDr?W#j�������B��&���ա���N�r�x�2�I�����^���o�4zs��wP9���/ ��vs�E;�חϪN4��$Y!�ҝ��O�����B'�d-�_-�u���#O\l�g˝��� ����e����f��C����0P�����.�Pe*�P�x�\����p��kpϤ;��3F��F
��>�����j��ά����?i�ޝ�x�?a	ǣAo*��5����V�߂�S��`ڨ��@z,����L�5�.������]R\�S�3�nU6X��+��!�a��̢�����*U��]�f7U!?��r����7�=O�A�Z��L&m_�����diN<�k��jMon��Q��!WË��	�C����P�0�Ia�(k
;b��Z�'H�S�`��q3�s'��Ee隸��K����{dWCi���Γ��l�k���|X�3���a;^~�F��_;�r?�Eg�#��̸巿�H�jN�mlնf����(8i4R��4v���?�yK2��D'� ]�?���R�!����o��~�|��ܐ���6��0�<�����X9%!{=�XB�|��_f���3g�D��n����|g�Ps�`j^�ɛ���U9l��^�q��yX&ɣ?�UJ����q}'�0"�I����x��mFŬ�Z�� �%�7L�<�&�\(1[�W��(s�l1<��8�����S���C�%S��c�S�@p.�ͫ�-'�(-a�q�Ё:���\Q��H��l�L�@i9�{��Nw'拊�Hz�����$|hF^�� ���'� ���8�^�1�Q�-�G�8fe��;B�W�W�q7 �n��!���ҁ(J�sWZ%��`|�����۔*����XH&�@ �����!�_��QM$�ܿ�;���z���W���e'��ľ��ʴԉ�w�h?��R:���D����C��x�:_��Zď����4�*�p�=�cH��;{g�.���.�(��WՐ�2t�,̺<R�f�'�dl�T���;t}=C�IS̈́�F�O�a��X0_s�u&�:-b�Oc��x�SQQ� �±fs��U�4���_�F��Ď��*Lg��+[;]5*�����uX�j%��Ӹ�F����̕�Q�$���__����6�������R�lW������^.�:�_ds9G�.�Eń��\�eA��84�k`΍�*�[;����'	��%��o3+��t����,"ӕW��Efk�W�nQ����s�6J i�)�k�DK��1ʑ�����l;�0
�s�F3 k�Dw#�ߠ�4y�Q�~���Ok��-��*4�I,d����lx%���R48����a���;r�
�<��V��Y�h-#h2?��$�u���p�Lui/��x�П�<���!�7����-�J����m�����֟e.����<�l�gR�?���(o&�p��D0R��=�A|V�:��~����Z5����Ww����b1�O���P�rk��q�U����{��P�9����Ι����ܳ�N}V��؄֯RhP�z�\��_��3C+��Y۽�2^U?z��X�K���">���AXBo�_�.��_C�v3D���QT ��b2 P����˞E2�oS;�
Wl��hSd�=��"�)�N`m�sg�L�SԮ�AS�>
\��T.$f�1pf�%���S�ѳҸw�R����&LF)�G��i`>�V�z�*��W��u�y<w.��迣��jغ�-I3<��M�O�g���� ��$ ��h���!ՙB����ɹ:���'.w �\��߃�t0O���sJ	r��Fg
5����K�V��.�f�Ͷ0tC�XBA��h� ��V�"9���0i��#����D�r��nc�0j.a��C�4��Cz_GϪ�*���B;wT��$��S��=w���["��޵���g��:yn#z8�G�L�<}�zZ����-5l�x�>�'ql"~�zp�'��J���x��پM��5/����Tg"��?�hwݭ�厩5'R�=m۬��ڤ;ޛE�,��m�Q#fҮ���iBz��v����j2
���+	��U�1��,X�����Y~�����y��ړ�њ{�K�/�=�;�G}5��	��.ͫ�9|Aj���$�i�Ȑ|��TWbe�W		�?V�/6񨷓���	��!r��kJ���"��O����*��`�B�F�:q����l��Q��q�-���sQW"��H8���Wװ���������� Z�Q��p
o�L���=�8���$zWݰA)2�a)���E\`Tk�饱�d>�D��GW�5Sp�ڪ��p0�C�����͂`��&���d����Ђ���p����;DFF��*��*��7�A��j/��mw��?����Ӕ.q{bZ�X�R�m8_v&�K����g4aC�P,yE��`g�m�]�ё�&����ut�:������+���Иvߖ �f��A�N��,w2��Oh]p��}D���T�����@�:�%�O����躭K�=����Tu�s�ڢL���0�����Tv�,j�8u^��P��� }��f��LI�����;u����C�#+�7��a��XB��Q.��d�����i�k�U�6o{�8����'i��"�𑭣T"���M2�|ߙ	/��՟��x2��w�\a��X��;�!������HD���_Ǚ���L����uC^��SU*��;�w]���E���%P���;�=�9
�v�q��=ct���f{�T�Z�e|�:�:d%�BW��|�%I�~bj�=|�����O ��?X>�L��9`���)vQ���(w )>׫��m�V����-�o��,r��5�o��"	'��A�Ht��Ϻ�RT���I�}���%��*�z1�Bg�h7٘?6�34"����ak	��2��2��8Wێ~��(+�/�fazvh��
