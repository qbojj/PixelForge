��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�06���A��E�T}�g_��i��WG���3v�gVO��ӯ'�6�_��őH	1h9�Q������牑��Α{�^Dߵ�YE���m�ķc����n	ao0��-r������)��rxΩ,0*�g��@[�Hl�F�/�7_&�E)�Q*]i�>9:�{m��X!�]���EM�����#�L����H@4������Ըc�3�HC��^������c&f���A�0���d.���`��,��sI�f6Ȝ<�A4�y���H����4O(��)�awN��U�2�3I��-��E|�o��{x��P� &��X���� ����{��aD2�Я����,p�5�Tp��SF��gV⎋��̙I����2��ٿI�̎���4��{Z������Bm"z��5k<�F�ܛâ�R��F�fH��ƨ���Př}�����b�� �ϻ�t�h���s��a����KS��7<!֗��@p&�<�aC�n��ȯ�XFn�*M2�d*D��Q:�8��y���6�wL��!I4�i�g��i]hSd��'"Q���#��ֺU���L�֑�K�"�K`�R��o��ye�^Yr�h�s>;p��n]�d���c�2�h~�V�gvÍ��{l V�<ú���9�?zJ��G�@_�����]HKc�Qp��&�O���}��iZ��te�U��׊;�� �=^��-�;D�?ޟk�ғי�R� �>�4����N�ҹ�h+m��  ���/wW����n����j��]�P˲i}[Y@�U��%��&zOc;�8 CpA
i�\8o������2w�r��Lk*�F�"[lz����ڰۢ�"����e�L�Ik��f
�S�Խw�]�Kn3���6��K�l��/���Y���*3���$/��X���#���rj}�.��<�f���E�l܅lٻ�t��e����lG9��:+�8�%=I���2Ԕ��R��5���t�g�@*d��Ս�z\	��&G�x[D��LR�b�T"�D
�m@_e��'�jUpWR����7P���![5q< ��Q+���P��,�1'l�E_��)	b��l:�s ���>�h_�po|�|��#d$��	aa���y��r�zk�6��u d���r�\ֵ?��١T��.���S��s>��I���k�ܤ��*�����k�� �6��H8�A�8��:]Q�O�@�"���׀J�[,��m�Q�Qu�{��9�| ��,�W�z�R?YcO�X������A]�T/�%�C������~Pu���4/�qߗ	r�����{:B�"�qR�@���k�����s���6Tz�cRlK�=����R�B0�q~/	TIQZx�t��A�ݢ��C���n\������dE^�(��Zpm'�Z�w�w"��<*I�=����JrCCG� ��k��5j���5�'��N�Q�;ޭ���ej�$�[����kJq�S��Z����]n7C�-Gq�2���yk��� ��V�p�kn3I���a�ޠ
�1�=v��`�O�f�Wl�	����Iz����肳�@a�X.�đ���Dj]n�N�>��S���4g�#h`�z���R��p���tS�5) �נ��S�����'��qu��!��!���"�oH�V���$�P�i	$�w�)���nA�QH�T"kƵ����{��H<�o)߹�P봮��3��,�����n�B���efNc�V˥�Z�a�w��Ղ��i*��A؎���֏	ouĨ��*����X���cD75�-�����ſi�Q������&���Kv�'�H��4F�*5֍\�z:���R\�,�I�Z1@.�)m&O;��U
��p���ŝ� ��w��Z��V�/:)DI��Ld1cъ�X��W��#�L��$M��w���V5>d�Cogurm��ީ)d��M��>�s��U�5y�_�F{�(��~�C�φLQ����L���t�H��ǖ�>�/�����u����f9[�<����<a�rkùT�ά��c���f�!�I����-=�*A����|��8��?A�/;k�SpA�:�R	�hp��ؚD��~�z����lX���;E�2��o��9��I]�KP@�,�+}V�q���8)<���
���h�Wb$�0�yέ��/|�U���$�%����Bo�R�ӷ�"(h�~�l23�e��������^q�����TN�n�@MM �pO��C���>*]���sz�q���^��S���-���u�i8^'Q*� �ke��fU���c��H�JQ�Ů%5�9��]����mx�k���;�H����p[�F��\�����ѝn�nߣF5M�^�PA�]v�3K��`��� �4n��z�ɳ�%LLz���fJF���7�˜J��O)A��}�)��nQ$��j)����f���d+�]'>�B�:V����o�v7�LI���P{��s�Z��}~�yXi�몡w�����04��]~�$g���Qd>/NJ�d�ͬ�"y�f]F��o�2�R^�3n�	<c��{E���"�J��$��i����r�V�mzV~?U�1KO��C�.�}�u/Ԑ a�G�����+�Mw�������+���+������}�'�ǝX�Z����ob :̊��'�xoF0x�Ǭre�"�k'nFyr�^4�T2�c�@�&�]��I�F
�FF}qrj�a^}�UG>���ATU�E����AQ�t���jA�k�0����梺1闚�,��H�ep[G�`<�:b�g#��~�gw��<Oԛ
