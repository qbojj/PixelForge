��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s������`\�3�*ME��!MܱO�3�{KIm��Iyn�C��(���JtC�nc���h��Z�?f���	s�qHz4d�ȹ�B���d�����.u�s��������<�Ś���O�?����b�>�[��Z�w��[����
Y|a'd�U�&z��lP�\_\aI9�@,a���60���n��v����t���(�V''�`�����JK��8�=��Vxci���[�Ԝ3��ٌ9�S�� g 
,_L���=�?n�wr�+���
K^�B������>����3�/��>��R�%:P� ���
���ϊG�%\�1���bع��2Y�&�kd���Ț�ÝA��Ɩ����u��ʊ�l�)QuOG�2j�y;�m���g\�f�3dȆ��Hq@.~����M}p-'�Fg�c	ފ������T���R�J��R�9H$wFb���C@��@��g�oA��������%<��u�wѰ�J�uΠ�=f��S+��<��*@E˼T���n��R^���׋F�%�-�x�$�/�W�^��uf�L�6�������V�1+ו��9��Z��VN?Xn�t��Q����P�j�$l?�7q��.�ׯ�~�RH���r<��ƑֱInnr�5lz����k�Uߕ�4B?ׇ҃��;�Ҋx�
�G\CS�=
~^T�X-,�љ�������ڥ�rO����f��pAH�T&�m�r?����ׄ�F��s�)�l��9��˞4$��Ÿo5%���ƥҺ[ǥ�ror��(���P^��4Gtc*��j�VA���^+	T}�ks`�c��y�/�e_�UC�z�����ʟ�7��G�Ay��+��7W�+a�Sv�2/�l���K0f$:na ��m�7ͯ��k[y�9�q���U�X/��'�Ya)�˓��mBښ��_�"O��8�2�y"�G�c*����X��,5�CcuF�Ȫ��#�0�ق4��CZx�9�ԅ�T��W�uEl�35��5����/F�U����E�%������3���k�OР���1�tD���S������C*)��'҄��,�B�;�G���`�Rݤ|����Щ�s����
�/NDN�dGY s���у}�Z_q�]��2�^<%�H��w�t�?�3�G\Q�U�|�	p�.^���˽�����&�]�C��Ć��({���2�M����T��z��:�j�Q(e�x�W��Wb$����G���˙�(|�������8�N0�3J�(i%�{�3d�x���@ݤ�B��p��	J8���Jˉ�,-�B��	��������̣��E�U��t�{�C�. �[�,�a���(Q%����^�5F��&'�zTΦ0�Z�D�^?�j/���B�I\b^���ヱoK����?� �~��r�/`U�Q)��BG���zLWt覘I�Mqu�����J���[	�5�QC!��(�@��-�_8�YM����A�ޯ����A�IwS
��*�L�w����e�����[eH�"�V����P�#Ο��S�Z�E�޿�!J��o�$A։,E�B��F�M�;+�nG#Fؓ/T�a��^����M]�X�U�a��K+'�Z��%)�ҝ �?<��~�"9qR���QX�|ߌ����J�Ȥ��_"w���/J�%�G*�q5*��s��P�f:�2̳F�|0I�\�:v�'i�Z����x#	΄)뤖�}[��M��.�I�%��Q�d��\�l��%+fr�[.� �<Z�����1�����F�2��R��8~*f��"T������˱=w*!#ϟ$U���P���>�1D�/��I�ӹ�B��ǲh.w�rΜ�z�1_*��J:`��� ��PF#�^a�O'd`���lي���L��3Z���,��E,��U"%����Y;� v�f���F�KӜ��6l4,��������kc���w���L��1\��(���O����D[@q�w�G�G���ã��q��Y��h|{i�j�mEu	6�j�Os�#�c<#�S�&�d��Cý߄8��I�kĹ���s��Xn`��u���,؊;��j�!94�`��e��u��xC�Ϣh��#?�$��/�RG�Z� _������r`{�L�,5΅{�%�]<lQ��+@Tƫ+�xysE>w����o��h�6[<&����Ė��[wk9u��!����5�����(���o��W�B��-�%	6 �G(1��]�(x%,HT�4<�n���Qg����XSt�J�/�b�5"x��(a�R���Q��Es��yۦ	�]9|rT8���
��E-]3�V�N�GﲧR-��?L������k���,�}&dTᗄ���:��D�6I���&����~z(^�2-M�Ȟ�8�{�B��t�Yj\hf�sXnBsW��(h���wP &�[-���q	����>�BG��4{�U��ǩ�
&�� z�,e���rK�n��̓��vm�������z2����p4_j��I�.6��Z-ݵߐ�2/�[X���X�-���X=̘;:��n��i�������(�K�d�L8���7kŀ4e7�l��Ϫ�zz^4��3t����J��zh��I��X��|Ŷ�6|�~�&��E7���7`�DS0�8��!,8����D�2���cׁ�BC�)��[�����X��a]x�\��]��\�;��ž�Q�/篮D�Zl�~�+L��:�M�E��\�����$/[|V[E	��G���r�rz��3�| ��_���c���gN!�>���( e��a����͉���h�Zte��@#�"��T�#��TS��zׅmy\Lq�8S���.�Zj�,�nb'�Vn=iׂ���}�͉=�8����'I`,���m�*ė�sbd"?u4�C 9��Hi?J�^Y�Z�&��i�:i���T0�ikp:|'�,�g����S7����,"L����ф��w(��O���s}/��3=�(�0����r���<߅��?�c^�oc)�̀�{y�yl�("y�Ψ�;����4�vj��ѤX�R�x��ȓ;H�k]?{f'�ܢ��x���c�w4�h��g��I?�=J�c@���tx�!��\L��n��0��f�����&J"�ǒ
qٜM���W5{E����f^8�	@�\������������sň�a&_+�6�-�U��c��*�D������1���� 5�9�1�xZ���׆q�5�}P���\�M��-�᪟�Z���Zqf�
��x�6Գ/���i=�#�|ũDH��2�s�E���ӟ6��;��3�bO�s��=��y����x����Ď�lu
rz��yx�Fܞ_^��^ƛ���g��j#� �%�Gp�9{�o�C�EGP����?"�fmT�H��u��
�ܼu}G��E
��W|O����Hjg���j�&ln�"0v����ȣ�WN�5�QU��by������Ύb���dеtfgn�YqN@yg��WU_tN�w��(-/�(f{���D�<O 5��q�tF�j�*�-����@9�Ey�H�xR-�`v-���M�bV��k�	,#�/�l�M�XQ>A�^L�[Tr���2�D&����K�=�9���aH}�*�����
���:�v�0K�����,�\zN�G���}#����y�Õ��z	FͤsO���,AT�0$��'����I; �gY�����r��BmiB�#�Ҫۂ��
����Z�J��*|�<�� �GF!�|@s�^�z�E���7h��雹Ԭ{zwC兠bϸU��.��!I����e������Ț�X���Ƃ�A�&��TDt�;b��/��Yqȍ���h�y�9<�����L��L����}� �_Y��*��n�N���d���"n/U+ǚ�	Kg�H)S�*��Q�@�XC��Ǌ�F ݾ�b��t*���p������߈wzmΙ�D;�b�ǲ���������-�p��p�rQ�fښ"p�W�ŀ�f�Wȇ���)�x��~�&Y�W�"(�|��;�dؕ�<�5U,�pB(���wۨ�l���n��IX�wv�H`�K��i<�T
���7��g�~ǧ{ڙ�xY�s�fb��F�58�K!*�7TX�0B������ ������ȳ��~q�S�G������j*� ��vݓ_n�,�x��;?�|hL�s��1��~i	���o ����ۿ*�I'��k�?�h��sy�Nk$�E������B��$X�W��b��h��|D�8�n6�F���=�I���+hgJ�;L6cz�CNxvȎ�$�@��O�	�+����qw���NS���^1dP+!sq�'�����~�[�i�d����.}#)靗Y�1�Nq�
W͈�?�+������[|��?�9�Y��d�;�+t�UJB'�[�/n�3���<"�k�a}�C�r߱M
�����d�psz�FP�$�mEZ�Y��Eh>��G	0.NB�#�m	�Z��[i��$�}s�		3о��m��%֌(�%EJ���4+�/�M��DJT�V2����u�"*���n�a=������%E��O��/?���6�X��7�ef��/�2�	/k_���J�p�UJ��.P���v����2���I�HnE&J6@"�"f���T���g�tӳ��M;��}����܁#�yiT�N"NFR�|��8��4~Ш�X�[s�"�|�e�E~��H�k����F���y�rZ�K�5���Oɪ/\Z,��?m�d���B�}U��4�;��^�:N�%�T�.�!����I��K�>�d��^,��H^,R��������+��[e�h�V�n���F�Ϸ1���Ҷu�M�ڵ�tD(��hI\R�oZq6Kp��S�����X�C����f���HT��F`�"���e),��Z��9ބf�o�3q!{�B�a�#ׂ�OWH<aQ��w��l��Az.�<`��oԌ��砻�P&;�
�����j:>��T��`>'	i0{�O����YQ(�~�>����L�g=B:ĸ�@���b��D/��e�p&��I��.uu��S��GM3scЗ��Żd'�^꺞�h�iN/3�Z�/��WG4�ާ�7>OfQ���\�*nmQI��G넜���Z��HaXF+�hc��Y�.�����⩆�����!^(F��0	����M��_��z�lؒx}�Z>C'c�*څ�7�mmu�>=����ߓ�O5E�ܘ{40�7$��oI#���'�7��у���:.���\�,e{	C�C^ B��(� =cen'l��}��ð���HxU���WB~
j�8f��,zp�H��>��|�����.ӗDUl�������O����j�Q��sf�c=[��_ž��~�W7I�Ȭ����%tb�cT�Zh��µTΒ�h���0u�Gӎ��/�qt.uj3�,�(�a-��6o5;��.O�:��g�P3 �i��g���C�� ~VA��i��9������川#�2֗�|Er��tp�[LKj0{�}Х�,g�h��~8�'I����0��9�� O�W�sX=eԝy6^�����.8�}1u}m�8�X�u0(op=�L)�ʥ����-i Q���vxkk��=A?)��+`�^���xv����!�[�L�D� E�v��,�[�2f-�����l�SԌ�$
px���[)}g�r�Y��=����� ��h><�>3%rx&^Q��������O:k��HOdq#�:�nf�F�G��N+$�%*�9L�VO�ӫa�!��#�D��pw[l��B�X�xS��t.��Ȏ��ד�A��?��a��{R=��7!c�}@U�y~]+Đ���o�L-L��w������qLڕ�{�~��6x]H #\u�иx�|{7Ȫ�!�$~�\~��g�>4�}=��o����@f��Z8�h���:�B���9�8���� $q�����p8X6�̍B���˾%����A�n���o�N:C�G��6����ً7}3=u��4c�Ne�-2���Y�6n��d�:؊?���ޔ���6@��7�ܒ�p��}LS[\V�G$e��QT&3�
��¤Yܵ���vB�Ȼ����9_)ג�{�W@[z���9�!C�/��m�$Sj)YnQ%+����^�Lg�0�1��;�
9��b͚X����6�lU%����&�ޛmSRn���[UY��9=Ѣ�CQ����y�>&�	��S`�#�F�>���.��R�n�A�j!>�a�N��|o[�3dn��C�C�_�((l@�H�b� *W���,Z�T"\��k�����U�E
G��4D��B�����`����i����֛KU�p"t��a`�j+�a�Ao���~��H[�ݝ6X�Bg|�L��<���*E�9,��!�E�#bՓ�d�H��'��wj�}:A(���.X�E�m���-M�1*4�֟�	�"�b{[WJoNl!b�-�8��-���7���ɪv����ǏR�2��m:9F�6�� ��a�]��=�g��5�>�����R��t{y�4U��U��Le������=W�eh������x7�\�����84���Mt��#p���VU0�]s�=ͱ{�T�=|�� wD7~�[��C�}Lؠ��?U��F|������-�����eV͵[�1�2�]ٕ��;S��T��p��1A0���-̮�1��D3]�-�n�m+|I��ߙ	W�І���rPg>�,R��%�!���Px������:�V��>5�#��ȗ;�0�UI_ِ��bϻ������~�r�7K��o�^A=EO��2;@��(��Y��Q:RpO<�P���I�Sc�3�ֲ&�x�M�}˫4-$ŰY;���'h���I�pܔ����W!�/m�J���� *��)�8�A
zB�݁�+z���&�g��RUA�>/?�;�e�G�#N�,.�~���_#��EAtov���o�b��~JG=̾-ʤ(���:��|���k �Ze�xţ�~/=Rɉ%��˯��}L�(~sx%Ee�x%��	�v�q���z��?h�(�|J ��>��<�+�M�LL|������j`���%Z@�uXSc:|�|��K�;5yx�h�<�~ngrī���I�g�ppd}\v����}=5� P@ϟ��?|S�	��,���+�%���W��GW��|�&�o6���SA\Q�	�"01W#R+�M5w���!�l�m.��av� �A������md/' t6�1[)���pl�ˇ�����\^ ᡾S�ѣOR�
�9���e�L	��|=-MT���ʘ)��1V�ׅ��7١gT���S%�/׺I>	;�n�ӤԆE���0Ȁ�A�Z�Y���t�����ԫ�Y/ -��+�D|�J1b�?$�/&����8��ߧ�I$��%�4��h�DFp`.t��_�Ms_szd�`�>�)��)��2�H����4�8@��+`;��W���l�M}(Wg�r����y*����,st�{��׿�-�M�e�6�#6H�I8]s�Z�_�j�o�S:�W���Ab�����������KkI5-���v�M��_�j&ǥ��(%��NG�	 mש^���^Ņ��:���s�$_��1���j����mFI5[%����0)J�Yg�C�0ʋ?P\�� �a�,n#�g�Ī�4��'Sj	�H�`VڑH{��q�A�	f����B�����H�kӑ~v%�����W�V)��q�_�تP�lcxnUgl��͖�*���1��o��3u~M(�s�%+�OT�#{��Ie��8�
����XC���Lj�j����k�z/�J����kX�f�篦������N��Ә��g�HR`n7��I?�z:���k&���=��jq�y�����&��dڢ"�<�	�Y;�n�R�܁����k��� �W��>��x5�t�l4b
OM������G�wS�Ka,�q'��^sA<J�_�J���'Q��	�CsԿD��ow��nN�;޷����,�O!����H��U�lb�*V:�=m
'"*��Em���a���1C!ȧ�2�8��UR#!�Ƀ]�>JJB&i��4R�[h$�B�D�gl(�Vk
��S�J��9Q��M�Čog��Z>�B,���+w&T;Z1�(HM�0���⋡�@B��O#؁�:d�7
J�)��vvF����u��4^h8	���h��#�;� 1}����$�k������8R��W@k*�.?.*P�,"/^���'�"0ᯃP��� �O����v/���_x�
���3�w��*�	���f|D1������f�Ԣ.$Q�"�5�h�����,�tA�g�p������сT����K�
Ņ�	�R�*�@�$�L%b���OʟE$a|%�O?$M���<�h�Nު��4p����Č��_i����/h����gEZY�AK�\_5��$*�J�Q���$+��y�B�1������i�|�DUI���q���t,�W� w�U��\qv��g�ӻ��G�[zo=.w	'rs�jAs d���"�
�l��B��ɦ��e��� O�][cY�V��̪\G�q�:~p�ȶN���^n������
ۏ���[P��g'�S��C3FꉮȢ���G�F�+CkR��Y���~"9!; t߯,A�H�/�B�;%�D���a�w��x�<,�I(��Xh�L���V���0'1�}��P\~�#�ExP7~Ϣ
�qo�6dM���b)��LU��.�9�MUB5m�O;�\��o��Ώ�ؒ�����2��H5Di���
i�g���4��|�X:�8b�)s=�K(i���5�A�8u�n�m""�ҋS�����t�l>��K�䤉@,��� �V7���2�����KN�q'5��, YR���\��C����,�7i�d��bG������PN�i:NVڨ���lVt��ݯU��b�Q�RX )jd�	z%�a� ��4��'�#F�P�
]��c��zݗ'�u������Ckf}~O6Ӻ��V�z��3������
�m�e�� K�,|�+�WdD-�:pGk�]�Ƹ1�==K4��B�`>�vQ����*�GJ#[%�Gr�uדtWU��gM�;��d"��R����?weV�������NBa^���w\�.�:?=����#w������P�3w|q����.�^���V��f��4��ҥk{��L�vl�~N����&U��0L���W�]��׾UX��s���l`\�/R�۱<�����xC���\��m�M&n�K��U:����kV�v��Akr�����qP�'����*�(Y5������gQJ�őc��qU�]o�&�&�u�����c6���)�Ez"E�{�
*:6�D����%d�$���G��*2�i�}ST}9��Q���2V������8ՙӬk�b@����Bڿ���qD�WҰ`�.^��r�8��	��-?�ͮ?ܴ�4ԍ�`1i&*"�>��%z�fi�d'��Czq�ȥ���輫�G-�|�B:ٽT&y|P��OQ2�X�&�׬�4ѻd����>SG�@^Q�C�N��$��������S�}�g� �՟*&����s�i'Go?��S��3������2�%�6t���/����(��/�)�`	��+/��<=���(�������b��_�b^~iZ���E�W�u�m/��(��0��d��n_8٧�/�����钇�~���Ѧ��I�`MJ`�*lUJ���Q��eCC9()&�~�'K�ɹ��N@����a53*�˻�b\��J��3R<�^L
�?��q�[0H�d1����e��ELs(����V����q�F�*m15��������=�7
}�'���JH�J�7��/֓Ŏ����栏St���}�Ɨ�t�~��V�P��7�W�e$�a�\��P �&�WA�w�|�a�x�d{h�E(*恹toQ���h&6�Q�\;�ȵ"�M�h?GA�����xž���6�L�ʳ�� F�%��uۑP�oe�� �$�SU��{��w��cq���b��*l���,{[���.�4���/.���kݠ�2@���*�H;C�M�qn4��16�0�y�~l#��	�-vr�Aw�M�A%�5O�@���O�蠎췐P�p[e�R��$eŐuv~L��M.��-<녘�x�,6m���lr�����X�Q��X�R����o��쉝
o݄	��]��Z����ɨ�aZ�ݛe�2��K��#D�;���k��������"��O-��d`MB�Ufa�z^ݒ�>�v|��D��t�ѥp�'�,���L,k��v׺X�^iyV6�u�"�:8ڟ�e���$����u���t��	�K�u#���b��Uǹ���D:[�%�a�7"6.�>����a���j��Ŀʵ��7�+M]Z�_��1�݉QI$w�1z&{���r��ݙc0���<�kd}>�6��(�\�����>�>��O�z��Q�ifXw4��,��X�,g�u�גS��Ҫ*����h�M���/Ӈ�}Yэo.�I��H��_��H�{і!)k� 	ܟt�$�7����1�#�#ձ��Ch�p%�:��V�j�Ws��F�t9� ���d�V�ؖ��vf�z�{E�����0e[@�[��2��3bK�<M�����l���{�>72���E��y�&h����)�JVؽTt�"����t�	*e����/�;.fڷo��!��S�`�k��T"�L�bP1�*h��g�ra�L1�����|sb�Š�
F��~�:EJH�Ȅ#�q�ͻ7�BP��w'^��}Q�P	�JfW=�D/^]]
��倕:�#��XbK�7�$2X��$F@��t�P�FDΡJ� �o�I}J����a�.����uta���k*�A�p�*�8x�1�� ��v� W�:^�� G�^��4Wzv��u|��v��-g�	�A/�	��>;�4H�~҇,�^�ר��S$��r�C��	�8�uv��^�s�塦��1��i�A,`��18�B2S,���\Y	۬iMZ��eBf�-U�� �`	Q?��^c��2�t�ݯ�9jRцÿe̐�\�Y��҂O��_k\��)s�l��$��H(�<8|��(q��Gs���O��0�[��lȠ!�<J�ۂ��m	�3�'��gj��H�晙:eh��2��2ץp��
By��V�E�p禺/�(����M��8�o��𕁏�R�\��(�~@<ڪ��m"��c|��5ZGx�{¹�4�)����v�`� ��U��]�����p��k3�m�L�q�.�Q	�����tV߁�%�k����l��'�;dq"�y�BI�38�9����i�7�uH��7����44�wٲ`p���r���u����ܘ6���$����R�إ��ٔ��?=쯰��.Q#��._C��-duث��B�ȧJ�1;���*�E������������`��Z����8:�l��3+l5DG��(�X5ƒf�N&�.Ӻ�U��4�? ���D	�h8�sCl��_����O�d�7V��>���W��;���DF��A�.��o��@�άgVZ3D�v�<	���?s�c796�	�ܗ�	����kNQ:��n�5�F��c�53u��h�Co:#2%N�яI�mp����`_֡<K�^�)ŏ�/�Hڿ���-���CGF�J�_DS����Y�̼I:H]���#����5~c�^�h_�b��A��a-x����4k㗛P��Ը�s���OGJ��e��|fY���܋7e%cZ����=�ڎGD����H ��0(� ����)&�����at��а����������J�St���B����]k�74T��h1���r���idq�f��a�O MX͜k�u����s�F'U�`Y�3tB�g�ϫ�.Ɓy��8nI�0cU���SK{%��!jv���I(2O��B�����͞�#P���K��q�����-�A��ӡ�hf,�V5d�/�:j�L>�b@/��/$���dg	���ĽV�/v�C"q/�blŹ�W)���y�}q�2"�7Y��ι�JZ}�N�A�E���ًr��G�����`��Z��%��-��9B�0\�~Y�	EX�o39A�-B$�!��(��<?Ȑv��W���DT8�v�m<5���_��]�9����>n�Of�giz�{��m�����ʫ�Oz0�w��sL.p,nA9�{�2���FZd�!l�b�eGt X�����ϟW!���-n͚r�"��L�Ⱔ��+�.���rߍKf���Jh���.uw"|���7}X�c����)�w'ʌ�O0�-.?I�:oU���߁�﵇�4S����@�c��a��
,�F���G3���P ��H��e$�J�&fG���+20O$޷OY=֦+k�pOA�+��]V*9p����BvTM�>{�I`ҍᦼ�1���(~֪1���wrh^&*^�N�}m)>��s��n�G
�s75�tF�������l����T����찈�Ø�aq���p�m_4@���
�N��"C#�=�V�@��DeH����F��qƞ����0�:V�d�cǡ��c�`p觲3���xbA�k�5���*����=�=*�����͟�ݞ��n��UM(`[�iȈ���um�pc�c���'�� ��p���r*�y��Q����k5E�<_�%�a��<1���R���ʒ��Ώ�D��ϡMeu0{UF6ڥ�*�y�.,�A��@��e9��Ht�}|����c��y����ZF_έ�{�_����KZ��on[>p��bo�\`G�IO�`�wGЁ���=�!`��/��;�Yu?u���T�5,�����(m|n��|�يԡ�9|�r��Go�W���o��*DU��4C��� ]q^*�Z�M��͒�����i.'^(����#K�P+��2�sA��^6�,�h	��j-s9F(Xl�I�{'�uXg�-��}�~�e�.g�?����>�N"_� \���cy��(g�D�՗��.��Rm)�c�J����Rd^�,�?�nun�}�/�����U�
������K�Wౄ�u���G�	p��ج�誣�pPVC�<Y�&y)�I�y�d*Jŀ�S\P�Uj��ۙ� ��O����W+|��WB������ʫ�������S]l����tL��Zԁ��@�D�Z��E},*���iH���-�:{�{k�r z�ވ�aB�qz��[��n�ȗ���@3mKa���5NXʟ��U�vB����Ϙ��Uû��1_�m�m���q�+�*{gb=�ڨ&S�=Y�����|_��<A�}̋ʷ�>��/�Oꗌ�HfXXwN��b�V)^�k�Fy�r�r�pq|���땙0�թ��\�Ji@=���=��`�au'�k�����4qt�hў�>�2�)~	�@�᳹��		��]�A� ʮ%r�޶ mƶ.����'�p
@��0�Ώe'ꆪF��^I	@e�
������s��NO+�H��U&S'����y��E�[�W!����&#��J��E^�$�u�O���CPAue���1����ϯeZ����6���,�9�`
��U�ŗ�y1�/i�2���q�r�Q�-���)�v	��@3�����5���h�B�0��5�&qx-�5ݟR�]B�/5���	�Ի�0�����!+�g|��C�1��FxO #?%K�v�.a�t=D*�Ъ�ѕ5*�����v�����^�> VY1ko�U�Mؤ�VGq��'jۄ�l3���U֜�� ���H��Dx�7�ݴ��t\�����oچ��	�~��$R��5��f(u��ظ���<�ƿ�^tmp��l"���,�)^�&�-��ᷴ�ϡ�/�W'���1����ϖ�z u����d��=|���s����sYC�W�x21���f(K���92W�j����!��z�6���G4=O�'�����g�ʔ��#���n03�O,�}����ӹuWgy��l�]��ˣ=>"8�f'�_"��Zx�����Ӛ�kTDl�Y�����0V�Y���M��f1���\V��m){g 6p���?������]h@6���P �Ѕ��������y$jbCeE�qM?��?b7�S�uwU,���D'ϹV��G���5\�Y���x��e~(��B������8�Q�x��w@.A��v?��$p��������oE�%�`�.\G�Qk�Z�Y��˚٩e�����Hf�^n0��>׶d5���,�P�d��L06�֛�A�����[J����!s͍9n�[�iT�C5'5���Q�<`"^��T�cj���_�^�D�%�7�F4�$野���Q냿���ꮉ���z6�z4����@�������|�������N�q(fa��h9�M�䙪�chN��c6���ɭ\�̮�⑚ҧٸD(��H��u�����٪;R�D�������E�ص���IL/t[��1Wt$A`��>C5�7�-�XS�^�/���y���7�Є����ß���!2v�X#���A�`vxd����^��R��0T�ϳ=}	�s��yE)$���%���x��yG���qj�������?���m��#F~��T���fw�S�ü������*�.��Xޒ)1���a��9�Mo؆��/�z��c%*�l�Eʯ���4�镑����*�o,2R�$��O���'�]� �p��������r�T��]?�oԸ�		t�C��Ap���p�=�{u�����{d1�U�HɆM�9��+O�VW,���i4b�,�c}2v״�0h�c���k��:@��l$4�2o�O�IHdA�ee��D��x�('>#��12s�v�_����F���%���|Ŷ��Th��`W���r���0A⾍�@Z C~y�����?�?]o�_h�8�����ۉ�����|�K+u�.o���YO��H��4R*]�?3�v}Cʲ]d�n:O4Rx&俛-�2>䈆b����MG�W���h ��Q�y���V$Sb}�������]`��lM��7�-]���w���Q$��T̥+7c'@\wЪ�w�H�����v�$L)W�����N�Y���uquƪ�PJ��մ���Ж|g��u���Þ� �BG)�n��I��҂-"O�3�ǹqBL*~q:j$:P��*O�1���d\����t���Jл�>/6�p>���q1� 2r�	��A���U�d�x��E����� U-Π��g��	��]�`��cq=sFO	����/�ouE>���w*��?��zt�����J0	�K3�P%1�l>�#K�_��j�L�m�a��B-e�0V���x�͛���]��(�!��hb�y�|j�����f�8�,FǢ�n&�l�xے��[�Ќl���jTv|&(H(��">7Q�T�μ�+�я-�(fFY|��Zc���ul=�q/p� ����&�az�����Ϋ9g���5�},����E�ȶG��"ϽP#�8�)�	NR�,��M)��"�r��3;ݧG��p��Z�(!��l�K�b�%2q��H-��[K���Ŀ����/,��VݶiWŏ��t�H��-:���[X�<LQ�_��wU(��$qU>*C8^4y�������_*��, 7�umy���`����D�\%�|�Q@����������}��(M
?/��}�F^���	�Kb�j�*	I���1�m����Ǧ:h�/j �_���f+�ZZ�r�8e�T0ˣ��'+��=��؃3f�[u��~DIG]����ˈ�n��"��Ɗ<��5�}�8��]�kzE��B�ܞ�&BP6y�>͓Y�GQ���h�O�[��S�@	����@q�Kn=S�ٲ՚d
F��n	�|Vcyu�x2���\�f����Z��I^�1�E%�kl��Yx��ytq	.����/,{n�	�[�F�St��\�S^�d�
���"�u�޻�s�13��Y�s%qA�J�F*�ن��ۀ�/��	h A��s|.��q��8p~#^m,q�˷�ާ��^J�� ���\�X@6�qD���E��ru��8�ʑBw��W��t=��1@=[ l���)�Y�j �0��M�ޣ���tb��Q�,m��. ʦ�ʰ�u��"D�, ��Y�������]+��aw��n�o/0/6ys}��l۵�Y��y�o4������	��Z�f���[��F�L�"7�<������/Y��~@��W(�R4*�M@��R&}�W���D(�(KS1��j��]kM��6 .�i�{W�f�h��5w�1"7�|�x�2��+��t6����Ay����|+�%=�"ﲽ���O�,��=��qBC��@oUG��X���7��}�n����2uz?���߱���.����¡1l�c��D�E�ֵD݄�)Bv��[^{S���r��k&:�(ȧ6�@vi�q]���#�J��"'P�`ۓ]�%�+�����.�a6����Q >�O^.3ݣ�oZ�T�7��X�F���w
܈�F�F���`7w�T��{N�:��[�w�+��Q��0�1�K�/�*#x���2�v܆#�U@�-���G��d*S�,��A�u����'T��C��b���6#JT�o�7u�F[%�e߸��\>O�G��Nw��&�bࢊAS1��G�X��B�1 �Yu�=χ���i�}v,f�]4��!}�=MeZ��� �
�ϸ_{m�~0˨�Py������1�pm(0�\�؏���P3,'~��n�$���~�Fſ�N���3̬�0���j�Ӷ�::�-{{8��2�@�N�z�����+7�/�&R�x�h(��ܹ����Jyоn ��7mnj0��x�郞�ӑ�Y�C��5�}	:�|��Q�'D"�s�����M��za�l���x}钌�@kV�L�f>r��rFՈnٵ�ת�X�`��۠�sc�4΢��|��'�ŧ9����+�c�t���:��Wl��G�D�,b�%����A�X&�'X���!�-�Y��e�S�J���� �,Q�T
�H柘�e@�X�͑�������P)���f�b�ԟ� X:���8(�~N�J")�$�pL��y
C��s���F72��[���5�T}�*ϲ�2�Hr�g	Jy��bCjL_�șM��;���E)F�1��Z��囹IdF�ij�R���cJV��F�yu��MCr<�|���8#1�}�!�Ɖk���A}�)��6m=7��@�<�x5��пxe��=D���~AE����L@��Q��*)\���f������dl��o�t&7�%�27�0�<h�#Q���cJ�^۱�=V��w}�����EҮ���V��+ҡ.~�|97�&�ۮ���Y�*_y4vMQ- �?n�P��Ê0�o#�PՇ������e���*F��:�� ����>~f����SM��~��D�Z�vn��� �o�zցd��u���c_�����H�AkM?�?��Y0A�ׯ���a�o�N�ET�_!��v2�(��Q�Bi�Nŝ87�,�k��;T��ɧ�����v��#LNy`�ˌ��: �tBA��4�(㏾Df�X�1 o�BFa��Q�s-���Π�|<'M\)�5.���"rf���H�D+�Ό)\ױ*Η܎HDo��P ��g�$ᵧ�u��9�'��yL*��#�@��`<��Wr������-_Ӷ���Kz�G��=�4���Z<f��\��Ђ��	S�~�X��+]a��ez?�:1Rd�����|�Q�s�'���D��������4^���Ψ�&N��qZ��[�3�T����"���ŤY @��>y�%��hI������=BTӯ/��=��~o���4�<.�:`�@�sh�2��H"�_V�Ӝ�|�[��x*�Qv��sW	d'�)ۏڎrpG�!����s�lW��������"DNh�ճK��[t�o��YJp�\<"g��ʸ �4�ѿFS�� s�mt�K�$o#�+Dh�C�f�VA�u�~�����4*;H�Jq�^����A#w�;V���D=��I~��6_��N<���ۦ�<v�6-���J����zW�����c3�7H"�gU�������w4<,ݑ^��+H����A���^,ZZ������vBO�0m&���f�c=��bV����r.����()as��D_�������l�M����a��[�N�`�M0R��V׻�Ϯ��`m�ʦÌƲ"��0��W)��g��Hɶ,�Co��@7l!����ј
V��u\����Ƞ�
�6��4JD1^�E	�P�p���[wOp��E���t��z������V�@�ЊW�,�O�co;�cfvV�_��-[��O�D x�7D�_��<��M�Ss�,2�੍�����f��W" 3昗k�4��I��V�4���� ���9<��[JM��7lƵՌ�)|	��B1i�O
��a������=��g7�9�/+��«a����R{;�1����7���^O&s ���6;��K~;lZ�8Λ��l�B S��ҶA�k4֦?�q45��?�]���55٥����S<u>0�$������l��a 
�MPN9��Z�c���;�E5a��ߟ�l�1�q$ Ӏ(��=�T&�tla���Mf��:�o9�u~����Z��v~)�8���A1��Yx����DT��lsl���eWN�=�ڄ�=��b�,�ݠ]���U��A�^m���?�!��jf��2z��S��r'6�n����^K4�~��*�p�^`��u;����H���<}\�[M���2m�T �gz�7΅��֧�
��Z���������9�������{i��8��'���oB͡�B'ECw�U��'�SG��x}
��l(q�'񹡠]W���W��E��T�f��ͤ^���X��v�5��?�0�����v�&�buh��$D�r�lC�	�)<O���EC>MXڙ�*��<��%�d�נpy��Z�i\p�{�1��������<+�&�&����V�c�P<EB��Hk�[pq@��)>Ǽ���Ox�)s�*D'9]ت��۠s�����PO3���K^�)������u��*���P�v9OA��N3����b,���!�1�U"�� W�V���g�m�x�W��O[�����B��������ѷ?&?���x�_�%n��a�auus�zy"G_��}6h)_�j��H0��z#���u�v�^�z�W��Sb(�����N3�w���D�99� M�=Y7 >��G'�x8hQT�L�L����#�-�p���|�x[��Qa{cgf=�$/J���s��I6?ۓ^A��j�ɢn�Dr���,$��uQ"��X�t�f�J,��0B���P�C��3�ֲّ��zv�|���j�nX<���lm�T@�l�o'��[�N}�Ύ�>u��NJp�Q�A<"t�l�#�H�k�PR� c�����/�TĴ�2�:j8A�Ks<�����d��7A�f��
K�m�tre���8uk;�|x�1o�֮H/�Eү��.͝��i�T�zu�}��ϖᚳIX�H4@/s���$�H� ��y:�9mn��Zx���:�l�m�G���eC���RZH8_��,d��;X�y�oP�h��;���I�Z�,"�� .�+$����m��b��䆈|�um`��xv�|����'F��{8���B��[s�a���x�1�VФ�ԛCFw�\���_�]�P��p�6Kf�+�[��m�7��Y[�F:c��Υ�>߽��N2��Kډ
ϦE*r�O��2n��K�lE�PFO����S�$	���%Bh�~��%(=�K�͊�QO˄'���Y>imO=S'B�:��D�2YVd�������������J'��
���J��N3Q ���N�!Ҍ��;�s�l����ݮs)��M�^�8F�[/��Z:��C���1{(B��(��G�''PQ���v�qE\
���u�.k�\�����Hs����\u[�8�`7zҼ����Թ�^�U�/EkHIۀ��T�͌>�F4�R�������fa��)���c���s�Np!*�1䣆&׉�2�h}LZ:�����n�O>~�g����0Į}�{�Ylt;9�(
v�2���1��4z%
�S|�+ĚH���Q���iN銊���~"�0��H����:������R��޹���M���s�g'B�`�a����|P-�a��~�q�q	�Z�נ�.q��Z��8C�6�Ne̗�?H��N�ʎ\fI�m����o��#�O�PS&�5���������w!3 ����v(��E@zu���9,q���@ڂ�@􉁋geXW�EɃ-8�@�:��Hx��YCm{̗k�V��!;��TP-w�cI�A��qjh��9�z�a-�ud�fV�Yt�o����4�ktK�_�/����30�m߫R fk��)�?'�HЬ���Ow���6�4�E�[^�I��9����T�!俘k�"F�쯠������̸*�N�2���}j�q��	{>�׺�}���i ��'QmA{s�[�M*kr�g#.�͟���K@�S0�Ŗ;W���%$����F��X��/��ֆ(�mX�؈BJ<��ؚ�@�����o�� �N)����Z��E�]���6�D�j��z�ѓx�h�L[������Do	��4�1�P���/U%�Y�Z5�}�)�Lr~^��R]�	ԾE Yd��.b���I����H��k�x���)�=��M����QŐ}���,����Sr{��څ��!#��Ds��`�fnܮA������d�*� oFa�T��!/�C��;�}^� ���ԅ�<fͭ�1I��W���<X(E����|sOwS�^l&,9p��0@�e��}��s)�����rx�e�="וr7.v;�M��(_�َf:���\.�5/y5���:L���8,�Q����.�\Ğg�w����1Tz��'p�w��9"�#�S���Kd�S'P��Ǎ�%x�L1�H8W�/)���;{2�~�U��������J{L�[��Z�M����ͳ}�� Fݹ�l�4|t�u!�Z�)J���?mr�a!�����3�.�^������$�-v��ʕ�髵,��:��U"�%���z�OL�[��GJ�3��y��C�?�pL|b��)�LN�Y��u��vŵM��:a�%�8��9�*,hygb\�t���
��^f����8���p�N�x?_C9`tN���y�c��]F�c)㬜/���� P�6��Q��z���+�"i.�2߱j�5b@�3�#�5��zR�n;�8ya�iE�΄:A�f��Z[�Uڪ������3� �;Y�~�Q��8�{O��N�`�	ؽ��f(��G���{��������?���d"���J�l�џ
�Nwi��D[P��pYz��u�����̮�pJ�<���Y�ˆ��ɂ,L��ܗ�sj.�{e4Yl�%諒�pK�|��R�C15ԷhVsж}�<����tEd��L�N�Y=�8Ւ։=K��5ނ�m=���J���Y�B�=��j�˖q�3�c��g��$+���ߒ�־l����i�:ްz����q$�F�D�.�sL�}��4��	�{>���ޝ��#R�F�[m�~�=Ed�;(���]\u{��J��6���v���K3���.t�9(Z\��e��{kp�Ժ,A� �)�0�D�[�HE�=�P��v���U3{�I�\����w�.	/K��6on�ܢqg�y�r&���.�(��O���]ٍ� .�#�T����r����x��Z�.�����1�)�ҒH�,���Ɦ��ݳ�%4f�wZFx�	�d7�:Pj5��c��D:H>�δO�}n��U.`�n�R�9X�l��/H�Y��U���N���m�b��<]�H�P�嵰���J�ź��
��]W ��y;B"��e;��i�.l*�S�F���o����'��o�C̄��ݲNt7S�}S) ��`L$;_�#$�Ｅ���]F�8��9�9;�	�CSm�G�m��:������"�mt��7?u��!�m�O�����˒�$&�s?|�2%/.-�A����$���f$0}�a��Z�mKD��g@����zvΐ#����Gf�ׯTeF��H�o%<�����������7>:�S�����j`#MЅ0�P���Ȏv2���^s���8.Frz?����pn{.	߯�&�*h��7����"P��1p';,v����8�*
��,��	@ߍ\���ݸ�x��V�
�E)~�w7VKʴ�b6l��'��+�I���t��ɛ�C�i��^�t�����T۪^;�S�" 麳䄄Ds,�ha\&̶Ӕ|/��+� NH�������8�,Z �H�SȞn�9�ł{K	�^
;��Nr�>4��a�U�6�
ֆ�lꭍ�Ӹ1�I[���{M���e�<��E��}���q�e7���0�d���C��|n�Ax��H4҆G����!�D��3�$iUt3s��ic��W�3�����_��Z��8F)]"��R�8)w�Ѻ僳z ��5
)�#�����d���!M�<�1|=A��!���x@�6�D,K:�T�!AO*� <�dx�G'5�.UlT���hˑE���W����U�6����th=CM�ڄ{�N���E�;YF�p�A�`�V����I��=��0K�+R�x�h
üF�Z��
�֥;"FT��sԯ�"z$|Y{�k����U���c����ܛ��JQ}$�w	�J%x~�t��X�ș�:���7_��t_����jϘf"X���js���8�p�����B%T>0>	e�[V�F9&^L�bٓ�Z�����zd|!`D�m�����>R
>6[G{^��; }Y��� Ϋ�H�O�8��ý?�As�KK���L���v�t	/)�n�[���q�X��=�f��6:s����B%�Rt^��w���m���(q���{���Pk���ۣ�Ua'�UF\6`�T3O?�L���)i���t��~}����<��$�9К���MM,zpuh-�\Z�}S����h�����p�n��XAW��)ҫكWU�$�Aŗe�̄N��9fN�lO����s��n��s»�!Oy#�'ƃ]NdY4za:����vĵ�d���_�J�2L��{�F//W[��Z� �dX�+���u�̷��z���NE���_�Y*���9�woV��i9pxL��_I �`*x.l�.��u5��iɅ.���T�-���S4 ���b�!8�6�o�?1�����B���0�n���{:UQf3je�,�C/�vKUmȪi|�e2@2�˳��$�T���}�<0���S�u�dw�ؾ#n�z�z^Af8Ǩ��� D�m���E4�ܾ4�������]w`8�D���� ���`H�-n�T��<ˍic�%��u֓|�m�-�X��?��i>"�o;,�(1�ۄv��`Z����SD�4
�ٳ,
��\���e��=�K��2�k[R����/}�]�c7?9Z#Φ�.��K�s�q�ԺƦ'��4��_� j�a�������@�U�N���nP�b�q=t�Z���G�RL�`��)A��'��K�C_*5��L}ဌzK�7�!����fc�{��{8��*s���wm���~�]��~�oU	��c�7E���s�"�n��E�P�cma&�Rᰵ U�L�iF󝯍v_�e1�ʽC�pR�}�������,��#X��mYL��m�Ҍw:���W.saU0Gy~�jZ����K!ϵ5��n/�a�L胙6��6e���"a[>�C�E�P��AOU*����e��A3LG�5 �����v��X�^ܘ0��u�!��� �u&7�1gK�h8a��i�"�\ih��h"B�gbf����F�M�U��IĸOf�u�R��Kp�qk�G���u����t�E��;L�_)��#b�U�$���|��^�~�W������jPd=8�B�g�ו#(�C�z�����~u��L-�x���фw�+$u3"}�3
˳mDO
�N9�\��s"���b��x���v:��7mEf����
ԅYvz�xzO��5��D�����?����3��$�}NNѧ<��d��a"G��^7F�]Uѿ7�'tK�v�� Yc��Ԣ��Z~E��(7����L�۪֤͘������"�l�'��T��N4z0�.��!;;�����ݼ����R=)~��>ѯ9[`)�J7?�
�^�:QC��=Wɇ�@�[W�n�y�9_��P����s^ -�v���m�����wc�u�Y���4����>e격��r@��H��!���@F��n�2+�-��lS��9ZӽQf5��ՠ�'�Mz�Ȯ���L�'gM��v{Z��y�@��:��o�z�00���c.|X�W�{Q��k꿸V>XrR������� 2�s�-��ڷ� �������c�@<?e%|��I�n�]��\8��Z��E>����b �5#���v��:8���#q��M��yUL�mƢ���Ξd��_����|�3owɂR6���fm����c��k���q�I�$��x�woc��o�P̩��k�Kꜹ��W��~������l{�#�hɸ�D��!|iHp���O�<���w������C �U��*�b�Q��p�~3�T�#IV���f�r�d�9�M��v��;6����e��x�}ҭ.Җ���Ab��!���#уI���X���x�'a[��F��	;Y/�&`f�E����b��g�P���S�����r\�W擖�ff�"-����� A
Ύ=��T��{W�������%�~T���/�M>�(�t�ZO7 Q| �vbP:�L�+'Ha�(y���B'^:¹wo)��t50�yI�ԥ���H�_0��xi���4Rw�o���%(��?�Tb/LI�Ѿ�Z}i����G`
���.It쵐[9Mr��nMD^X������xU�&��O�VX� ��KxL?�TZ�H\H���1�d��h۪7P�����wt;fY��`�%��fFJ^Y[�>��Q��d��q��^ݖe��~�n�D-C��Luf���"��N��+�hYw�t� ϧ5I�f����D3<Q�_,y�nq}z8�7E�=j�ӎ�x�����egcL� V���n*�=�)H��ď���! �~��a��^���>;�nEw���߉�l�#!rg�n"~�Sǌ�w��>����*��C!R�$��J��8� I���:�c'����^E+,;��Ж�s�]d٠�Db�{�&(����F�0��Q�ʳ��+�U6"J���֥[�T�!7�Ր,�F�6AkU�\��?Xa� >�#�+h��3�'�(0�ᤧ띉�3��C��ʿ�E��K_9Q�k��x�l���M`u�ԫ̟��DG��(��N�l：�%N0�T�c�w_�*����JUPZ��G��ʆ����H��b��Z|9�N�k�E����:gP�b�$:�̵�?��{̃}�R(`�s�=�&�2%��҈�4dj�g�~��o�m��d̊-�~��tǌq�ڶ��������a�ʈ��4X�}6�A�"+ ���%���n��O�y�O�毷���[z�(����<Ӑ��Ƒo 9+8��՚�\��A^۠�{Fa
���Fn��Ր��
|�e����� �[��b�-����F8���[����++�i���6�<a���1�m�A�:(��q�u�`�K���qK��5�Oo�5��䧢�_J�|<��o��ɓ�Y�22C��M����.l���t	�+7�2�Y8����ږ��@�_d�4q*$� @M;{���F�kZC�+Ӕ��=��6�%=�� ���6�P׋��p����1����t��GU���d,�$.
�>_z�bgMc�fo
�௺�U��@�պk����g��"�R��5#�n��8:�� ���3cQI�_>(��ԭǤ��JZ����NYGkI��Kӻ�uQg[�c�a(��O�*C��U�0Ŵ��$��.+{���qu��ի��q��u��,��0!u~���:���䡲��V!v~���+��}u�CZı��A �##�-D^����d��ϴ�����:�a3����yK}�hb|��x�M��R�<	2�� =X��Ϧ�`)3�M7�p��xpSw%4�j�뮲΋�8�6��k4��W��=�>'�e%gǓ@��+G���-�@���c=�}�Ǔy$�f��mmcI�D��22��֡[G�x��׎gB��oJ&蘭�9P)�dl>���;/�V�2�ct����a�KH�#UA2�@s:3͑mqg�B�]��@�/-�B'�Ue3�{��ؼV,i��4X�-Jʐ����@4�җ��#��w O�G3�o)�����4���r,�Gy?���6�R8T0�k�EgS�#6н���+�Oi'ϊ��]]���Ș��(<kӤwC�M����gμ�V��lu�]JX�������O�sc�id���\��793}��q۝�$�u3�['c
