��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��I��i}6�_��Rf3&q%0��-��/3B|��P��Ɏ0wk�N�Fy�p����u ������cS���ԸV�z;4kƮ˴V�:���]8j
�,�YğPѾ!����M�E��������eg�RV���_w��f,i4	�����0p�Lܧ%}��떁-C�F(��~�ޙ�����~�F��-H�¨�vd����n(����v����6��/̇���ҮƐ�wt�)w�K���;�K��JP����
���~̔�b ����h�]�kGtub���&���h��5{��n����CەQ����� EM�T�����H�?B�/^�Ӗ�'N�
�K���#�.9�C�x��\f�~,�)F��|)m�u�_F�X�gÃ
��"7y��-V��c�o��o����w2Zi���S[N.?a`�[7q� ���N�Z�G��X�u��	���
���mx?a��x�O��j 6$/�v_�{VaL; �i�WH�CGl�2�R�W6U��P����$�c����ߒ�6�B�¡3���m����f��b��1]��V�G*�j>�a0��������f�u:�Ҝj��-�l�n�so��{Q��T�N���"{�m�*���� ���6����/�^�X�_�Q|R۪�&V$y��fR8 %Q'p�U�A>j�a�Cb�	AOt��RZ2��J�ӵ�G�g�DX��7�ch3w�$Di���Խ����I�C9�3�w�k,��3�$+KJ�v��|u~�2���ʭ�+u�������9�q��B�$�-}XL�+�j�S4�w�I�cͤ�G<F<�"�ݪ��0Ei܄�ɑ�U���ts�	�/"��D�������������0�k��|砷(�g]�I˪���z�J�%Sx3d��=,���*[h��{������;�K�j�����Ql�"r��n��¢�[o�������!,��˵1B��i2��`�klU�P��{��ܟD��N�.����L����2�1~�s�����g��<��
����E]�����tp,͘/�y��6�����9mYۛ�xU8�t��0v�i�M�~��8��_D���>�� �cC�w�)�΋m�.(G[Xc1�w`�po[�6릍g�zW�Ɔ�y T�h���W�Oó�Ѱ춒�`�﫧���4&V}�����^��VV$E�.!�e0`�FhNH�d�B����t.���Gv)<yj��3��;��*���Bz6�$��FZ��e<�+K�����"���i2�J,�3k6M���D­�}��/��n��4<%�O�n������� {��~��(� "��9�[��J�#P�4���6������u�e���������`��\�R*4��EӼTӆ���q�����|Yo��cߎ�{�Æc����=vA��O?��V+��N��������(�g:I���ݛ}�`���J���=�7\$g����Qoʊ�'�1����t_k�4�r�:b�؂�w�s�m��5�KE��X"�SL?�V�G�$K�dcG�������������&�Ta>+v5©�a!�Ц0P�o�$+�]p�{�Z� �tWa�NȒ҆9�'���q�\W>�dwn�����(Y��R�F�W��H�Q�M�lI���GC��A�O�����V��_��7�:�*fs�&7y��Ս;}V���l��1�s��@��$�����f���¯m�V L� �tX�������q���h���fh�X��z�i�(AB)�Ĕ�������Մ1��ߙ�.��7��O�1�	z!���9���I_;��t��a<�>NL��ʧ���� �)�S��9-o�s(��Zj��Ӫ��[���lì�n/��@c�%��m����?1���ɡ���`�=�M�Ssru�r4�(f
^��}sP̢�#A�
�)�y2��IR��� ��^��/���+�'7W���_��'Z�T�(�&H��~Y�ĭp��b�?<1��&�������2�)�}uqu�]�q1���+���`"�(8o'�#?��!�aRa�㲽��}�"��x걒waQ�n�g���D�_�.̗��9]?BD��=KBRzկ%�3}���y-5B��m 1�K�,�xl�hr�x�xZ5	N���PFxSZ~��>r����gߝ�W�K��xQpg+n�4��\|r�B�c}z-��2Òd:�d.]f�\�j�I'����jC)��sl��<HkE��	��OqJ
�}w즰��l�R�}B�@������p*,��կ�HJ��:CH$5Mo��Ph@��_�����Uk�F�,<U����LC)�Ĉ���=Y���Tz�JB��S����!h/�z�u��-ޯaҚl���I�^��b�E�i=��"�$�2�	1���|K(��r�gϻ��Yc%�n7	�������R]l�ڠ�d��c�|(�f�9Nz���*��V���],&� 
i��!p+���4�Sd ,9]��K&x3f�߂���q�������X�/��<�,�I���AXW��4-�̯>��Wj�\�Ӂ�l�j��'p��j�K�R�v�e;+V���2N�-��4yv���	�]E��D�/=N�@vLI i��5��/��'��
v�2��=��z񉶓X�:��y?�xd���O�O��v��Qԉ&����q�D�����c����;��u���כ���v��L�>H �5w���s�:� Z�a�0��� �Gѻ���V��>m�ݺ��!�]	���R~�ڃ�?C�R�^���Z�cԩk���젡_O+U�Y���t��B�j}{l��uB��?	��ӌ,�+��������s����!@~_���H��7��Z�!e�v�i/�oX��9��X��8��e�,�<��v#��'�&�z.��Μ>�%�����:��w��Ư�zs�w��滥#�QB��`�E�9�r2r0tʻ�в��,Ѥ�a�E�D7_��w��&�Q����K�9�����i*`��|�:GT�f�j	�ZC湠�liz:F/%�$��Veq�r��۱���Ec�6[+�~D�z��1wu)��NS��W	���)e�`qE�?ӻ��)�D�T�H�V��������}��e�<j}b�m�uM���Q�����|WF�Mヮ��ײ	)����i�=/8`\���eQ�>k�h��;)����t�2$d���+�zr�<�e��X�4¡I�gf�v�-��us�{GEE9����A�"�ƽ�K�H�\C�,I!�Rdy���I�������BR�z��~���G�0�ͱ��� �cT-�c ����貽&	��6Zm����H2!
����?� �1=��a��X������XFX�"��K�������'sv'Ŗjڙx��c��]>q֕���yq64��˱)�����Dz߄`�&�ld�W$�.�E�,�W�0b���ĝ��<7��]�m�������/	 �]���LO�����l&yB�/l�8�n�w�R��OM0�I3Q�8J��N����+�`���9,��r��u���L+�w�ĕ4Z:�z�sxu�
!D�{��E�"�	h#�k: h���a���
��i}���ha���Q֤��e������h99P'���B\;(N1�(A�d��zYR�x��z/B���K�����7�5�
��`���H���x"{�I�@�VW�,՝K���B�2��w|��w�n�nH7;7?�Q3�p��-"1��".&9��N��k�6�p�G��c���0ǻ݆�|��:��&M��l7�����jq0ec�nX���N��z��ti���}��
�[-�V�ק����E"��@ݻ��~,� ���:LP����X5�h��}�R|/.��R͛��g5���x×����<H�n��5�)�&\��%<�g�$Lڮ�in���bCVM���&ș�l�RE���0�&�s��k:<���ߗI�j�p���^>"�Q�+�
�ښ(�{����gw�`L
`I��Ǵ�Y�a��r�	<fKO}������ց8E���`����QW �A�D �"}�/��z�f?�`X��}�<�H��"i�m�3�pN���rf'�w�L����|�[���Ue����)k/�8�D�s�ݟ��T_�p�����-�~K*Q�Lk�ќ'���ȥ���f͙�
M�5�9�ekn������}XX8��r�Y��?8k�I��$�o��9�TL� �r�����K������n���/叀�#s�7�_&��DC��Z½D|?hL����fd��, �ya�L�TW��̓"�_��*ȴ�6QגK�D�%�����m�n�6e2;1�f>���TI�RG@��c����61�' �����YS��H��{��o	�l�����0�t ����Q��������D�����A�I}`%���1D��:{��y+h��[��0:��UYs�'��D��4	���|$���c��+k�!���L=t�����H�ZK9��mzV)�5���	b����ȁZ��oI��K,4,�,��g���rL�y�X{�Tή`Z�F�L='�G���`�2�p�+�isT>�@9�y�B���1��Q��3-�=Z��I0�uE�e�Ǘ�F��k.��D;Tz�{�R3�yOC�
�2|�`��fW��$8��g`�^x�\w��"js��O��ݖXѿg�ȝ�oZ(
5�g���f��9#�f�0�($���WY����;QS	��!�kn�N�۾,m �s�c���i��֒��M��� }_�17Xw���/�;�J��"�j�I�l�Ǿ^&H�T@}��ݥ[�B�5ꡅ��_5�=����nvUF_MDp�!���M�Ug�2<r�����d�ow�+qb�|��m���Q)isޞ^�ӑj��=!6��} #Y4�p$+����&2�ݑ�� ��G�߸�1�l�yC�sl*�M00��>���5'_T#�&��7���S:�e(N7�	� Y��@��z�P�1꽑c{�1�'(;�&�iхqA�3U���d>�F�>(#H���G	�Cu�y��(3�Q�ݵ�������:i鉞x��wg����b�o� L�P!ќ��V˷	��0I��P#��gO8�;8�`�M"%y��|7��=k�,����V7{�����#�5�s���|^ܷ1}Q��N�VS<�6$	�Ն���5���H���S�Td���@]=���㐷:�s(x���o+��vM�����0���]h�,s��Uz�V�M��1\���ٰ�~���/�a�˔8��o	������Y�:��Z�+h�UH���NK�h����3y#�J��,��&�̄��v��N��\z����15"��Y�����4����Cu@T�=���	뜨�!O�,pP�D��j����.�f4iՈ���xS�b����Q^VDJ��S�֪�݃���_z��Ok-$����cR��%$�����㞎K�7jL��8c�q&r�7��b��Q��Db���j7o���0�	��_��\�
������	�$j �n�( +�eڕn�b !1-����T �m1��K!;�$�C�C� X�F���
(�W�+���U�Uc2j�~m6����t Yǹ�
,��m�(}y�͔\��r,ȫD/�渙=?ƳQ{�? [��
ڢ�����D/ܿ�=\p�̱�֎��,yG�ezU�08Ll�o��#��Yv����[�V���|x�ۀ n���Ǫ=��@m��.:+��d0��l��w�x��?A�	Z�;�%;Ź3���%M��ܣߠ��*}��������yk<L�����-QH� GgL����n���<_�v/݃����ܱ��׍�I��U4{J����*G�=��@;�
�����u�K�
mB:�Q����2�l YkMiν�vpA�r��?js�5�S���`\�.M�����)t��<�
�����q���S'�f`G�݋q�t���6zXH�C����_
�XWB�瀄�g�����0[�H�e�,��rZ��b�e3��~so�[��=�9���Y -ק��Ab\����Co�P�φ�26��9f�KY�ֱ{���4����D��\���Mxs�bL�ͤ[��YM��Axf#9��K8s�K��19>f��a�Ch���a�ە��j{���v^�Un�c���#���ɪމ�����M��$G}І��2N��ϛ�G��B�(��H�@�MYw��#?����-$x�[�.B��v,�2V��?�Go 8��7o��@&��&3�~������GtA8ס�q/�R?�X������<e2<?��
i��GdF��r����"jpq��<ع�wQe�Va����F#-�y꣟α��ѿ�d��͂)8�׍�K썧A��Ԟ�ڑcJ��^��nOƩ��$°9]
�����b�.���������L���Y?�����Á�����S�7ɍ�Ƈ�ٯ���tæQ��?;+�V�1�*e�u��G��6��^�"A�zs�F�RR���>��Qɗ��^$�����8T�#%	��t����l�P��&p�[�U�G�|��W���7;�X��a":�V?�	f��
�}"G��J;u��viӢ^��g��p�%-��j���Jk��3Vr�p+sM�w|�Ȕ4v��ΎN#)be(��˳3/�qN�����z�J����]�!�<D�RQU,?���7��&W
~���aR`&�h����Ϛ"sJ�_���O�r�?���p�D�II��}��
k��jj����'��'�Ix�K�'���6����Fߊڻ���e@B�ٯ��mp�p��$+���Y�E�� ��ɫ���� �̈́7�P��P��[<�I�O��4���
�%�R��^��T����rv�+�k��+����y��Ǵ��dT����1�@!�<x)�=�hTAV�k�O��Ug��ͧ�b�t���A��E/�YX�Y
\yhE����U"�����9�u F���.;�Sj
q,�������oS�4�G�3���O-�3�F�������K��LD��F&=b�la�K9`?�*O��\��o������!P��a2Mn'㐯�Ux��i�2�R��bۄ��C������1�n"�`�H��X� ���f���$�&��2�v�i��6e��_x7Bğc�;�a��	a,�v�OGO���S��y\�`}�ؖL}nT�nI�<��K��؏�S�b��סo-������ܟ%�koIK�P��kF���KG��y*����'nh'��1+��Kv���)�/P:rJ�H�����UQ�Di����Vڮ���]\ba�r��&)gq��4ԨQpo<�ba<GB�NY�=�L�~����"�T멞��7�x ����2�',�I`ox� ,LӽN�^:��`)S�4��JXމ�M�!�ْgE�B����lN2h3ISZ��G�F1J.� ��i���N�s0^,�;�L)�c�4V|����7�?����G�}��B8�އ#�s=���ȩ*1zN8iQ`�~���wX^��SC�*��o�Ow��!�)1�C�K��ai��Y��1*/p�NP��>cϦ�Z_H
:o��c�D�V9��h�.M�^���-�9��`�Ş«B��]��r(s�I�v�G���i��.�h$�_��}��!F� �	���*B��SP
�+F1>��o�h���d\r���((��̖�$��x�2�%��\z"yf��l�f���o+V��m@�v���%��5��\s9Uz0B����a�d���!��_�C��!��A��iF@�_X'��e]��T����z�k�X�\�<j����[p�paA2��&����E�S{�c����|��]���,���x��*�u�)���M02[%1��������3�t�=���ˁC�H%;�#�+ݩ��w��i�����"����o��јӖ-v���kC�^�ڥ���<(��.��o�(�r?����T��}�C�C���y�pc��P�t6�Gqg������U	F{�>��@�C��ξs+O���p�Q�^�ݠU�F/ϏӇ�2je�c����Zl<���ōT��#@W]�!b�)��(����6�&U���W=�y �B,��]�M�@`<E;�6��vx�ZR�S-Y	/\9K_x'�J �29!l��F���$���ܤj�!�|�΄�U�E��{HR/wE��<�
?���ך�����f��&��B%cZy�U9��3�H�~��; (�W�hY�a���0�J���P���@�JI/���c���!�R~?+:]hZX�J<UzՒ���a+���&cQ�Jo�4Y|�F���1Ͼ�e�F���1��K�������,��W$���qa�5�7���t��RT���ow}����wYc{4�ȯ�w~���s�HQ}��D]ThL"�B&h����+�T��F�F����]DF:׸a�kEd���1t ��'����a����yF�r�-"����a�>�*׳ȇ��?H����qf\^�1{�a*�w�)��Y���	Ǝ'�Uc��z�����I�|r���%U�+���_(�+��G}<���'�ع���9�����r�n�m���ΗUS
�-#
2L�Q�0�-Xo�i�<P��8�%�ܴ��M9�B����}5s����E�Qj� ˖��wB�Y�1����RC����C0G�6Q��A�[�����ˊ�Z���Ae[��������D��{�nA�����!��9��k��îEW%'��łgbl�~�i��
=@�o�vc'gm��hP�1���ִL��t�=5T��Rb��O2$p .��:-�+�yp��4SA��/�'81/G �l�q���呞 H�G8A�:�zb�Ôb�@�����V��
(�������T��x��r�5�
�[)'���6i
N�!���X�P�<Ul�U;BV���w]M��w�Ǹ��H���Y�>8��	<n1ULGe�������st4z��u$G�(~���11���FG�l��!��QrJ"�I
�	����������O��ٰ:jà�G̽<��b�ף��b���K��
9:�{,�g� 5hM����� D	8nJڻqW}~�S��5rTW�+5��E��GqD�v|2u�hɅi+>g�����m���M��hj{
�%x�����\tC�5<o�l]c���eɶ[���ʴS|����x��}*������
�x�FB�D�O4 %|��j���pڐ�ެew��O�R��)�!D���~���w
�Gu����|�ig#���L�
Yt���e3s��U.ǫ (5A\�������~����٬ԇ�����HW
���z�z�v���H=��{ԿvF���♯<��ҳ�ү�z��D���Zݢ�h\q�߆.����Wl�g �͐�=���<
^ڴ��"���[|�6�Ƴ��M�a@n:"yT�����8��¹Ţa{�A�*�R�R{�	3�/��~`�J,H
u�S�'�M��iX��v�m;[��L�ɖ}Ҝ�� ooG�z������\��)�W���<"g��,U7y�@{kR��_80����V3���ծI��Ծo�������(���u-�VP,��T�Ō��W�D���=�qp@�9Q|9���`���c����B ��#c�A�P��*v���%��e۝o�|�K*���p�T~Ƥ�_l:�L�� ���hHO'{pǤ���	����7�F�b�L�pjD����W
�>ej�P�j� �|�(�{41z�l�X]�T�[���m`Y�[�a�+����������WL�:V}�I]��g�c0�sc3���[^~7T���_���ɑ�I�
�/�W���0S6sD��8�)>)�	�yIe��Y����!p�c
4%�DF|W�*a
7ߝW7ݛ��c���)�s^��@B�7�K�<����d�#p=]r�G`�9YN�y�k1�6�h�JI���7�!�����xAfS�Cl�m�F�ֺ!|�j�EK�����D=�j'\��k��(�N�c�3������M���%�=��	�~���l�L���L�1����,@�W��� T�� �)��梿��;�m���Ib�N24�(D���zh���n�n�Ȯ�� 	6A��Q'�~�����.���;�5��¦@���#T��Ŵ^��IP/2�3H��:[�t ��P��<i�{u�3�0��r�s'�k��U'Ⱦ@�*(.�Y�3�xg�=}&AR�� ��\�>)2L�S��G�ťKd�!��������k���Xtdg�x�wJ(�+%��\�4pl N�nWS�:!>^Yr~d���g�9p�/�z�����<�03WB�xV�K�
ac�@�V`#�5Ju|u�l%�2.��1w�4hњb�-x6�m �W�Qr��Ъ��1[�!��d&|�g�/2L�x����eC�1f�Z#��̮�5y��n�����u
��/ %�BJ6Kpvas��S����&�ևv�G�V�#�1me��E�k���ñzv� �(��!�в��L�2y�֨�&��u�#O�\uϒ��������m��]�N�Tϔ�݂�;?��x�+��F-��(�}����G�FOVy��V@����1�v買���Amn����G�G+A8+mN%j of �I��Q���p-�j�/㔯��J��� z.�
��T�V�iH�dk���� �w!�j��!�[+:"a��<DH"&�\�G#�;�XĲ��О�ؚ��=��= �̝?�����j"� "U���p)��G�ǱU��=���3RA�)�E
��VL�!��M��ÍB9 V9C�ҏc�c��s|��+g��c�C��ڵ�~���ԍcQ;��F[Δ��I�|�zQn ��O����_<�[|�GL�"&m�R�(�8&��Z~̔�lN#)4�W�ݙ�]�3z���
