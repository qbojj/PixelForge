��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0}@���?s����H*O:=�@�eQ���-?`�w�GK���gJZ�ݔoZ%1��s�;q��O����e��Z	_����h~�n,�ȍ?��.���c����R,CEע���R����� �A�<`�ʅ�8Q�"ױ}��T+:C��*w�En@�Lj�k�O`mW�ԡT��0���α|�Y��M]um��@��W�O�j���2b_0P��6t'��ϦJL�}�#�,��|�w��Xv�v������Υ��b�wZ|{��^�UX�R��H�[K>�f���R��Fֽ�C �6Pr6n������^���a8�R�{�3&��o��-�5��ҁ ���FTfG�����ou�4(_(KDZef�z�V�3�˝M�O��_�U�KDwZ�\�X��m�~�7�@\J�oM�������mE���LM.~��KP��u(Ĩ5�&P$�����zlW��𫾱����1��7D:�(d�;�]��=�w���J#�Va�ۄ����!e�
Q�z�M�����N��SM8�ga����2�K�/�aP��l�H1n2_s�C�WǇ}�ie�-��z���1ɼn�n�e���K�&��
)	yU���:�*|����|�p+�0g���Fq����l𨾁�6�w����O�j��5�R��މ����M�h_lq�]q��E��CQ�#|d4ڹr��<SsQ�x}֌��T�7�����
�>:=ď|�(�$M�j�ش�8)�������@���T:��]��)�!�x��YiM*N�۸��xp��F�2�~��d��-�7�T�l.7�3wi�r���r�u>�;e;Dw�]uK>U�p ����g�����g8PPg�y%������"6:��_ď����U��|��+j�lQ<���x�"�3!��;�����>���;Ӣ<��=h.2�oj���2uzV�&oS�B��=�r'k!�/�Y��� OyD���=�Ģ9}w ��na�Hk2��?��9O����&���N@�lͨ�C ����f�i�I��z݇޷��,�J됯Ľ|�����U�r9x��6�t/��\��Q�l���(����RmH���j�}!��}%��Y\h���֠������\Ij�����L�$��P=�D�(�� �_��rت��V�PS~�9��4c�+
=�%����9-��~P��ݣ��ƏvQ�b����?O�,��2R�?Tr��A+��2o�6�Y+�\�`ťiP�Sj{E��<�i�&�S�g��ۚ�a�q4J�;]�����{��P�Ͷ�TX���Z��`S��bT������3Ѣ�E��Q��lߒ����F������>`�<�����褙��^)�}R��7r��Msa6ǒ�d!�|J���8�ts�I5����:l��IDY�|�Y5r*�b,��>�E�I�~�=�9_!Ȕ��J��ϱ�p���C��F����k���Zl���W��G�6�T���P�5 i��1�2�1o��8<�[v�;�B��͜B�[v��5��G�?)m�guiz���-�G�����I��룦 3VAFE�V)���UJ6�fF�I�7�[�t�`1���n�1#ɰ��t���]���u\���#���t��,�Z�UY��0xӳB����i��eS%�|&����N|�Xr������˙�* }��L�@fc�$P�t��&+Ҟ��R�BO�gq4/���uI�x�m�"�Mӷ��Cy���: 0����)^A}ڊ�u㳵#/��Cٌ$7��g��rj�Ȼ䉉(�1�-���B�bZ+���G�ri4��)�� �_&rm��J����:�4����>���-�+�0=pp�!�q$8�m�k�f�]tVo��wwr-봽Hx
�/�'��|s���s�U�ڎBٱ�9���#��	e~>��%�_8^�� y_�G�O��t>��_���E ���]E-	�ƛ�:ǻ�G�㧞Z�-�L� \��u�ϴ�u�r�4�G�&����YJue�؋�-�Zt�3CL�;�◎7�wj/ծH��'I��~-A,Kj�Dw�
�+]�@h�U��N7&��h��Y��*-Ŝ���9TOV��˵R�cV�Z���y�_�䴥<��x�l���j������3�F�Al�2�������`LkW:����g�A�ñ*�PE:�����P�u�ԑ�Z�(3���b�<��dS(ug�+�?Þ���KOg9�V��Kн2�
