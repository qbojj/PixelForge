��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��g��C�$	�Y>|�Q;^_ޢ�O�_=W�Z��V4ST>�.�z��>��� �:�J�/�c0�O)4=qߡt���>G+O�G�$ $x�6�=�Yg�Y<U�t�T#O�@���{��7q)Y,��H���f�$F���Y�a"fM_ ��<>+x��1�:�������?�5T\������z♂ѐ|�b��T^$>$*��I��>G�"�2�t�O�wws�iP$	��l��&y��˰%��R�oTБ���D���c �P�L�O7�'��\1�t3��4���c�A���t�D?#��I���ru;N|��M�eu�+ъ��Sp��(�Z&H�a] +���}I7m�5L�n��&+ץ�D�G
$����!�=���6�I����R��2{�l҃�E��E[B������_G�;3kI}�Y{��~C��{%6fqN�}��L�Ɨ�~U?�\q�O�o���$asZ�3�Sׯ���7��s7奠��6T� ?5Қ��,��F!u���lII���X{ب,�];
a�u ̧#vGy���%�"�
p�I�/��=��,v&z��(_��C�r���po:�d��0�OLܸ�l��I&g�;�"���g��V^������S���(hU�Pɪ�Q�q:)d�nPԆ�����i�I��4,�59��lm_����s5~���8LDtp�z��.$L��ҾS5PA�`L�G���K*�Q� �>X�4G�9�}�OuͰEa��FeM|�վ#�����9��0=\62EZ"�%��֖��!Ơ	�PY��72(�W<��I��m�C⡶?�S�J\�J��]�	���<�2}ւ��]����w��2�T��^cD����\[�nn)2+��}-��'���?�L��>y�P��$�AC��t�Z�/���������eH��pǩ�1N�7�J�ʓXUVb}��'��w��Mdol�J�;�4�������n��N5li��в�t �39�?cع����5����$}#���թ�W���'gOG�[%�j*`��+�<ܖ��4	B�+��������Ҟݲ3mN%$�0�D��x�������no��qde3l�ݖ�f^ z���H:�q��/���������zG�����dS�����F��N�_s�j��E#'ΰ�Η�
�`�X����X�B��C��7aLɤ�r0jb6�&���j e�k�PcXa�楈M(#U�tS�g�	�t�%�H���6�I�J$חW��Q�*�Arj^��1[�=����[�٬�%n���l�K�(��?��A�o�{U�P���?g�cD�|G¯�~�JR��c[�w����	ȯ�e���H	����s�2����
�a�p��tI����rO?�e�a��I+��6Iڵ&I�]\+�rܼ$�?π�?"���:M��ɕ�6�u�U��F��{@yZ_if��֦&�(t@��;C�a=�Yh�Ŭ7�,;�d0b�D�>Q�I�٤qC����4P�����!Z�BD�a��O[�d!|�gD��u~������ ���t���k�6GL�n���^��+g։Qc�O9����j�9��h��w1oW�)�vث7���H�a��g�?��|r1��7������G)��fi�8��G)�hՋ����>�G('v�%��B���+~�&�|"�*W1��X���=����$6���ӨNj��*N�=ć�򩘜�^J&{�v�Dm84g�h��Iv�\L��Zˉ�&kk��V���oJ�_\i_�m�r�P`nH`�/呙�%)lO��$�~~k�H��W�8m�3����q�d/�R�Z&O'�\�"��E�����̈��F
e)o����Jw�ts�t/�y�P��X�����Mf�r�X����;��lɲo�*83��8�u~/MȊPa���N|(��JA���8 zN)�%�I����[��N��3*l���=���1YJl������N�p#��j�3������������#]S�d	�jU�@ƿ+���>RhД1	F&+��ƐG#�<�%��7z�t�N>�I�˫�')�0��
#����:����r�w�d���b�w�܆�DA�:�a��S�F��?�aU~��
��K�$��9��P$]`�]�Mf�:r�sІ��_�{�"�:z��Q��ot
�u� <��VJ�=��&ηh��Wץ�T�d�k�a��7�(�����Tfzc��o����`�q����8���9=�2��������<�Vn$��R1��_$�Kl(f-ۈ9`Ϲ �M{�j��ࣻT3��>8y~�����a��K3���|��iB&e@���4}H`>��W�Ĵ���ti���H� �������4�`�z�~�׃g~�����^��F\r���C�H{�7�^���C�s�Ͷ�#��h B���,��r�;9�j�'�kt9�1"��wS�j
9$�E��͖�Y_8�Jx�a�j�)��e���خ�h���(�u@��I�W��q�����_~�#�� ����8	�t����e��@FR�j��7�A>x�p9�c�)��_�eN�4*K�d��k+�O~biT��E=ʕ�<U��T"�2x�C���>�e�}�Νm��0����� X��0[_���t�=��bk�������HAV���Ay�)����|�� ��m$�e*�ċ�\�L8�;��1�%	��}��6[��rP�b��q�Ϲ3��4C�s�f�"v=�����f�k�\�jB8sw�N)$I�)iS��5��&w�D��v��= �ɩXݚP��x,�N�vg����WVct�2��=։@�2N���݇--1$�dZ
��foP�H�Ȍ侹層z>��'�~:�;ފީ�(ָ��:�_�]�q��cm��/qp��b[��N��G�|����TS�u!����2۲>q7�F��{h�c��!���0	�r��}�+���<�`�I�4.%�ڂB�N�<���~�|	�!Mk��H~'o��W�2/�r��uqRH�G[��Of��NE������wDN�� �e��(q�PLD;�6o��
�1| ����i"7^���,Х薲#D�m�R��=L!ôkpdn�$�d+B��E��Ù�� �$��]�HFzA��o�\�;a��;%�%����G]��B�@_�tM�ZЈ(D�)܏�/;�(E	O�%�5��hAu���w0&�S��R���&6��|ol���s&�Q���]��j�=���^x��g�H��2���:�p��@�%�R3���"�3[X�t �nHX��������1kt>���<�n0��&ȥ� ����v���s�o
��A���ċ}�������(T��`. ��}J�9_?M'H�Y���Y�� ��}�Z�0E�Q��%�hk��#P����84��sɥ�v��E$���mE1�*^��e�,w��I9�P���P	������O)�t^I����u�����[x�Q=卅���6Y���Nr�]���E�w�돱��O���\�HCD��x^�LOx��r���$��Dw7�K�E'�䖩��=�Nrp©�r�#�z �'x���ӵ��;[A0��>宠"ZgȞ�l�Rn�]���=���]�q�Ǆ�Y�M��p�50ӹ9����@�9I���G[N(�{G�P�)W�7��L��{�j7�H=1��	�G�k��$D����+�'�3Fɑ��I � ]rÖ�2hA4FU]���P�fb�
iW#Y�_��j۝9yII���ܮ�`��c��d��J����◖$s5j�8��|7&�������;yF`jfV<��h�/6�s���Aԫ2h"J���O�L��0���udX<�U4��Q�T���w̺6���R�r����8�!Yl5"m��aecC����hk���&!���p>��x�x�r�#��ɯ��'�k�$+���n�vC�y�~�:�Հ]�:5����wj�XxcKS���;�zT��#���o�F=qĳm�j@L��=�����p�䭏<��>]d4�0�.R�D�c�<���j�Q���bbT�ox�{��b���0ye�bk4iv7]x`hgn} ��}�1(Ij��'��u(?t���bx�O�h	���(AVL� ����T#�� �V�/'+X��IBk��ﷄxa��d�
�w�Z����Q��Q��iD���B�t�n�ma��J�H�s���Q9���� ^��k�?���C2�.]���?3�c�kTկ�;��O&y#���F�%Fi/?æ�4���]���x��A,��\�rl���=��&}HzVcHMY%��VǠ���4lfO���2�&���t�Ѫ��O�H��:�?�l3�y��׺�$_����3۪���4�����ta��j���q�uTH.�_H�h��������	4
�pi!I�A�:�Y�n��W�<T�V��[zAT� X��ly�T��W�*�]�����������R3/� ��d,b�����$ܪlyr2��dXy՛
R����Z��Eu��U��&L>ڦ�|�
FdL\�X�]�	x�%��"uu��ז��o�@���ݗ�5�#:�a]VI~�nZ�Zz!͖-]��fCKV�7ݱӍ����l�e������Sד^nQ��$���Ovw�4�י~g0JW�*�����G X\V���w;�(L�[�F>�#��7�^��hH.v.'f��J��aW&�H�M��Z�*UJ.�&?�]��GGVt  }%Z&#o�F��#�8�>�]\u��X��΢����D�LE"�x��-��?#u!�CP���?���z��{p-�;�l�����@�s A ��j�%t"[ҷ��ritԿԦ�:	g��Ȕ��e�4���U�[����i��(�ٲ��@k XB�s��4��*���?�ͣ(���;l�*Og9߷�Η♐�BSf3�>���?(��|@ܿ	�>u����BM�u����M��Ğ�L�|��5C�W:]FK.�~HI�l��%q�1���Qm}�B�,_cCM*q�+`6x�{!�u]����G�:�w�)��$h���M�����S��;��KѩιTڲ��c����P~qb�4�2�1c����C�@;:�ҐL�}��7�lZ3
��X�*>���(�;�c��<.?zJÌ���fâ�h�	z�����'`#��>8�o\ۇd�:�0�@k����w|)��Q�����'����l|~R��k�\�����;ɍ�N˖
���z��!6D��sQ�_S�s;um|�jC��D%��4��H(>f&'U�E�8��d���4�b�ͥ���oX� SF)�� 5ڿo��ͨ�J���c���H*�:��/�j�T��d!N���내��d_`�'*�n�Q���S�$9��W���zP�C��x?$�~��k
���;��>��pr$ �l��z�u�#<r~��(yj⌦n�"�b�6�fs��ݔ��l��QQ��`l�f���P�{��������߱ay�N�V��)˹�8���t�E �?��^l~����h�J���7��1CO��
�tr8���.gl�`��3��=}�@#!�LH��}~�'����(��jc!������������6�#!?����@�AV�/%yO
�4]+��.�b���8��k��{|�|��mvː%r��oF"SES�0�p� 5ĥ��q30���E۠�0�p�ٺGt��`��g�o5^=]���rj7r ;�<��R��؊�l��77c��Y�b���}>����3�v*��X��$F,��9��'��Ⱦ��C��E�\5m��#�����2�爁b�	�V�|g�lM
���Y[���e����kk�F���?�
�:��|�$I���h��� �GP��4��B�h�'ù���РZhբr�W�v�T\�I������ц��荊=t>'e�	F����s�	P~�I�~|^���J��?e|��,#�W�_��T�z�/������.�Xj�N�;��)����ܶWu��ϡ���_m����=��ܬ��ckӊ���U#�`��VJ��p�����HWH?E0'��m�3�c��J	��"8)up;>x	-�H��v��y/���ݮ���c�2�����bC4VkT���n����`�k�I"ŉ/���!��e1�q�|E5a*:u��u�a�;\P�>���jIU��+�uE� ֊�^zú�K�����0�U���BSA��XLǫ��t��/�` yoo��U��vm1,W��`o�^���Y��`��4G.��	�]`�_}˨��|Y����h#�����0RT�,�윁kK� Nw�ˆ�0Ƀz���>�n65N\s�o��p��cL�#�.153䕼�)O~ş�������n�X:�Fh�V��Q��a�W�*�\@u�6�;��U�7q|o�>����>0x�P�Ϯ};����
�ü�@'؍qY~aw,a�y�zm.�y̯�s���@aSZ����C��7~�"29��([���5��ȱb�9�q�kdq+��L�~�\����.D`��A'��X{_���ߒ&n�3�uxC�x7��%�,'�$K�������� �������+�ٵ�x9H��9�k|��sfF�(9��g�Aǭ!�9�t��(�8/[��KK���?��i���-t�9�i���,^��s�=~uU�����[�B%X0����S�Fu�Yp�D�4��`N���Aכ������t$��d��3L�����ฟ�o������!�}�'B|G'.�����ܘѷ���.��ɓ��%ݗ��N��t��?z��1	��`qSC����(l�F���D	�y�2�퉇��S�:��>Q����C�R-��~A��t���ă̵g���9�ۘ�e�X���t���z�jbf9�>Fε.�Ç��d_�2�|e��/��Hֿ%;�L�Ӽc�2�JW{y|zs�b�X7�N�WR������F�T�?�;��>e�TT�<���I�x�	��X��.y�Tj̛��]�d�F/�#s�h��ux�A�'H0�X�AZ�9)W!�$X� %������J��W���AI˵�G��H_�A�j��u�N;���\{E'�6��@\�e�l�\���`o�cf��B�E��3�@���<��멍��W��@"���U�c�^�����jo倫������cL�N�99��{�ϒ�S�*��RQ��	�� ���~�zӓ��������X0��|M�+��|�{�� r}dv��}�+�q�=�O��£�e��;'�'��0�2��hP�H���J����'L���Rݘ,="�えl��Jnc��s�U̷+mS�NgB[j˶@���LϹP	�|�;�܉�9D3nv(c���&�h9i���m��PQ��Ul�pI�����;w�ضz�Z�>�Q���d~���Ǌ�������iD��*Z�v�X) <�AsO��L�j�KH�3�5���ܳ�����At\�ߤ7SO���?�!�휕D� �����&�a�C	�sD/p?�u��K��گ��f�D�>������sB���>xn����x3?��%� 1	�u��2ՂQ^��j��j tg�TL6D������0d�>�c=�%ؖj3+��*��.l୪�ͧ�:��c���X�4��D*��a9I!�x��x.��ZS*<�X�)��hb�
)�Q���]���]�0���zj�w�G2���@��)W*E�㇩���e���ר��9%�<�;}�!�Z(�Չ���cb�k_�s��B̳�=������ �hmuyBo�uR�;k8E<개�}�G~�yf<��1WTH��ޑ�--��*.(�bhHu�_ro�݋A��$<�6��Y�qH��p�>�=��b°ۭc���cS{���͗��=^DC�`���~9'��=>����9R �J��e����c�+���'�)Pt}8$�����J�HVI�hKw��lv�G�C#P���޴_!=�n�U��{v�' �K�r����HV��I$�7.����+��R��]��M*�����!/��@"��\��vj�e�2�_��x) a�*@b^̏��9
y��\n�R[�@�Z�-4�A�^����@Lme�u�Ap	fF(g�]�1VSn��5$��u�0���8�V��"ޣ`�f��[�K��![#h���m,[A7�5 ��+�K�C7EO�Ȅ(k���	d��ͼVi�tK��ƃ���K�9a�A^�e
��	��?''�Ǟ᝔�9k.���>����Y�W\���G:N<\Cbv��'9��9�W��(vr}���S�x��3���ٲhj?+x���ae�������˥6�?,�ɪ�X5�(M2n��iJ�'���T���>�;κ�������N|�����"F.6+�j��Tf&	��k���D]PDs�ZJͺ{����*<Z�^���q3�����y���76� �ʯP>J�af��hͶ"NRzB�xܣ؀2��\�w�X�Ͳ� �Xh&sCJ���;��ˊ$_H8�`��w%<H�J�`��Qi�	�3� �DoD5�x'9���&��2�z����;,�P�;]��V���Y�&��3��ݑZ��`֨��;���lm����t���J��U1��pf�wrB���B�����i)��@�h��� �HL�8N(����׻���;��{�ڶ?Jzj����`��g_�V�35�گ#d{�x�L�!�G9'
%T^�K]�1\�Ob���X&���`��%O�Q��H%�?� $?a^uxL͢��T�UB��o�(�ק5��H�B��x����k����"�xPe鑟h`����ș���g��d�ڡ��?��:&��r�!��-@�7����83�K�oF��{7h;��F�^6`3���P��u돁���Vs�r2��`HA�_�%B3����f�0�Pd���7e����[�HYƣ}�M=B�w���P��=Ƶ�J�(ʩ�p��@��+@-\���lՑWv �#���iAFn� ���@�E_�=��� ���ްe���.�D��o])S+f�J�����Z��b��{v��Oy����d���"$]c�q;�%ŕ�Eyj�>�m%ڭH{��\�. \�q������0�Wy'I�;E�wո�q��$�� .���mG|� M�R3�ʐ����&�Lf��ҧpQH��hs��2�'�i& ��<��1���ג�,n�܁��]j�n�d� ��3!�}[N�G
�N�<	a���9`e�������Ӭ�=�x����؜�ܻ$$hI�J5޹�'���8;8���J4��u��SyV��G��
�A;���x�F��@Ղ_)&�Q���y����\ݒ�Ʋū����YT�q#�&���V6�����\Uh�Y��b�$i�H��ii3�������x��0�6aP�^�G'!yB���W�;�v����R������!.��^|QB�pL��ZW)-i�ZT�����DC��R����1=��S���R�����+CY�ȴ	w��H[����epngT�E�$��>~{wTÍV���Q�Nt.�x���ќ�.ʭ璆�+�Kn�iڤB;�H���P{��~TiyGŚ6 Y�}�����:q�1���.���ٶ�A:��sdN�8'������'��՟K[C����8�u&KEuSw�@~��ȷӉ��8X��l�>\�]�F�gd��-���$ R�Κ�R<���H:�|����A��!��'z{��J3% �"��yrO�G�w���)	D�i�}�Χ�>�e���S+o�ڠ��W�U>3��j��$#�I:��U[� ���ΙB�1a�J˦`v�(�r��j�?�WXs�����㫂a�=>�0���<�X�=TX�7��Pc�l_������CC�W��ܝڲl�OH��[��,ǆ��.�H���]ll��:Y���?�z�(Cm������زC�ODX*Z�f��6�:�GQGВ@mV�	��o��A_C���r#f5?ϓ�4���d}�v4�H��/^���X��)��U���~���ZKf��Nv��~11� �7݇�]���ծ���p�9$����M1���l��V{��e�9	'7����o�Vǋ�&��ilW6_�X!�$��-��Q��{���P�3��CZ�ym"�у!�G���Ļ8P�������&�_�s�� @�D�%2���l����%���@���rw�.�PHT��֡H-���)8-��:�0��Xᎁ�m�m���T�47����w �/I	�C�,��\�F�j㷙! ;�ќ���w���կY���ρ�P����1
vLB�3 w�=
���EO�����O��!
����)�<�b;4��'����$��u��Kj��-�kU�-?���kpD�3�(����D���rS3_��Gt�}ǫ��$}�ZbXƚ%"����\_D��-1P��6�M1|~���b]�+����!Q�(m�%��X�L����۵n�X�Uy1b(��*v^�jK0@nQ�b�$�߅�R1��8�h`�+Y�h�5��vr�E٦��{ ;.�T����Uc��&ق�"�-t�`�TC=뢶&�>�D�����|g����)��_ۡ��91���~� =lHe��6���2/Y��Jl���	5c���s"A��a7�O5&��&�:�"�)�3F����Ed_�����,����7� �E��	�g���!�*nH�q�|�zmHΰ=e��,�Wrf�5��4tH�G��jC�C��7e�̺z�[X�T�걡��;�zV�#����� 3�7�q��'lu'���Eٟ�of֥��r���H�ی�@�p��K�ռ!{�)^�k!�0
b���1�eH6�<£��4�d!љ���B�[�2lw��ɲG��n�z��e�{N��\�A����"-��M������)s��""2���\X;E37*�KKQ����Cط�S�+x���F�XA�շu��C�����:D���GN]a��dT'�����-�O�)(EZ����?(��S�X-ރ��Uk`r9�yb�yf9��V��j�H���qLH,�»�{5�ݿ2����ZDs$���e^b��M*�BZ ��o�Zz�)i*��'�����X�\�>سBAe�W�b���j$�6�hG��"#�APh��)�
\@���>+٥�P���擑N6���t�-]�O�:fL1k�:�{�_k%���`�*�e�x�b�O!���d�p]~�b=�{,��In ����^pe�)΃im�0]�`b0��vM��KaЉ��2+�]� ���|�|]�T��5G��-�ht1�(��1���K�-�&�g��F��8��\�R��ѓ*�k�,��Il�F��	��W��I�\����[�=ۮ?���/ "_P���jk>����5�v���;)(gH�!g/���*=����`�A��Z��i�^r��S蟠Ǔ_@��ˍ�poJ��>�Ћ���ٷHp���#���� 	DږV�����<�'N�U�� 2|ƣs�(.긋�[�D}�i�~�nL�Ow�>���#-R2cHH��'wܬ�u��3)�i�.��O)XS���R�
JA%Q��|�)�3�i<[lW ,�fz_ɠP�QR���5���6]T������T{��WL̰��m~����T݀�;�;�F���:��/3��IK�lg`c��u��+���?�X�B!�I[RY��9Z�G�w����-<�?�o��ᩓ �Om�G���ȥ�T�hf`)��pi��/fP����PJU��v�?]x���a�X�� d��4g�����h���M���D�e���P@Q{[��4����w�?Am�2�[,�ڹ�\�����l����h��šE��$�L]�|�ʾ���׾��&E2��ei��cu+�jw��W[��
�}��yHl��ܐqϷ��٦�|�˃\��۱8t˴�q��M�(� �?D�a��ɛ���J�z�a�K��]?�8<QQao���\�y�M���#$�u��,�����t�`�h!������2�?��`S���%����ѕ=�ͦ�4�ܫW��B	�B����hE�J7�`玐�p�Z�����şla��z|ē]�i�78��7���|�䯷�*}vv�E���δLW}��^�hpf�~qkNۉ�f^�qp{V�A��H��6�^S�"�����'��^���WdN��⤸��� J	�#�]��cm�=F&�,�!]r?��.5���@��ׇ?c6���k��N5~�:HX�I!�a��c���ixjx���$.z�H��B��et,D��m�uv���-́��'���O\��(bN��F��:z�eś�����↱\ �T����+&Ih(=�S@1&�3���Iy]�R�v�t��˔�����a:����9�v=�ˉ�|� ��}Y̞{��В�5z����ϩ��јx"A(;�$n���V�w�87����#�`v�}+�Zj������	�V����� �wX��R���k�m�3N�|���@��D)�&�=-;�u��0�:���	_#%�+eg�@s+6�{)t���܂Sʌ5���"�Ւ��hă}�OZ	�dP���m5�3�&��E��ٺ�I` �c�������v���b����xbqB�b��QQe�{�HG�N�lO6�f����k|�]�����d�φ�xe@)a�ũH�;]<�*�
A	����0��)zqf����#�0��u�'@�w�np��,�Btn����.=G���5􂁿fw�~	b��#邺즜ȸ<T�|L��B�1��Z�����#���o.!A#G*;�w �r��M=u����e�t߶�]]�h��C9�tp�\N*rm�r�'5�Q :i`v���G���x�������#��n��|��']2��K�S�ٞnʂ�(	pC��>���p���*q�PL��VN�R��ӓ���
�*ak"�h��R�p�
�����1��6F��l�,�OZ���b����<9�et"�rS �|�l��_�֟v+W O4��P�J��q
��I����}斤tp����q+�_Ck�+f��tnr"h��4��\�#�������:����Җ�[��{��wJ:ts$�U�F��6�Ȟ[;aq��3�+�z���;�S���1���o	ZA�Sݷ�w���W{�1�LXCw�
�;M7�Ʒ���g%���D��B�=���
B�@M%���`xQ��pEkR��EQ�}2u�=�%,+։��h�?��)QO˱��|:���EJ���N�뺌䔫��
)�������r���FeJ5D���72�G�~�>ڲ�7e1�$p����5��^�ihS�r��H�<��*�KPð��>�2�I�c��xナ�M�w��=�	��m>���*�J�lN+*E�N�Z�j����F���7��j��x�ǽ@�Z��aK ����ؒp/$�ޑ�.�����&���S��*Aӆ�1\z�wW��$?lJ.��u�u�ݽ�-��Ga=�| R<~r���3���'{Z� R�Y����z�g��ë|.[�Bd���$?��~ޝDO@��I%h��:�`8��b��F��Ċ�w�Z*=��a��C�#3J(.Q���u��H�0��Q<����G���)|T`�SɃ����.��l���2��w�i��gV�̞Qa"����:�0����������t	~�靮��y����ÚI�i��P�`l<�:�� ���yKJ=���an��tP[D�M����}����\�S�����â�@h���*��<MĊ�+�*F���'|�?r�m}Zc��5tg/���^~ԫ�LN��/������I*�52�	�����a�F���;U�����\���,;(�F��xף=��jz$R����c�K+2�"�L�с�򢜸)J��Fx���L�R�O��̰7!a������:Wv9i��?+�����ӷ���$�@@���0=���؀�/��T*�eKlǡ���J���_��E�X/��Wsf���hR%ȵ�N�GZmQo\�y��f����z�R��]��nk�>�hX�N�ySU�;܌��\\��iD�t?4 �xWYn\Q�K9���Pۊ��c?��v,��]�*밿�M���CU�BX�l�s�r��D�R���r��F*�t��2�XNd����m� 
��G�b���|L<�͝��NH]�z�CT�{F\g�Ev����+p�W����A����Ť�_A&Y6��Y�0���o���Pf)ߓ�_��0�Lc�p�{w��a�Ea(�Vp��u������̝6Gi�9|x����fLlg�;Y�]� u��Άf���=����_��N[L�@�K�CJ��t\�(�a�l�5F
����\'1~���N��,*���M�+�.Ldu����OИI-O�����'��C[�4+�A0��������J!�҂��v�=�5���4�;���^I�	�ԛB��������b��p��`[��8~KX��ON���_��:��Qj��p�Q�M�Ps�����$�1��&, ����[��g�n���D�	��У�S^ /�n�OT�L XA���v���X��8p2��#�`���I�0�����L?g+=>w@	uǔVM���#	�PΗ���2W�X_�4��y��7fA/�fd�E���`�XY^`
g��{��L"��=/��|����CcU�ab��5��=�'� M�9Bʼ�S��OC�λ+�m�-W�l�����.�k#�*�R��L5�ji&�w�ݷ(���R�Lc�X� "[�O8�7�r�լ�-�[Z���dW)�Q�&C��4�5wd���Lň�RT���u/l�N�M���I��#!*��Y���8�(�E�n<|Y9�Qt�`5R6¤�I��m�o�7a���r�k{��(�y�I��	E�yu|J,�3&̄�w�X�2���/�v#J��� �I��G�=o��u�LwaB����j�h�(u������V*�z��G�x��V'�֚�	��sگ�X�Ž��q}�Q��k�A���q�nc��#
�~|4�+��Qs��j�m<* �(�hA*uW`�|X-mt���12'�]ɼ�UhŹ&Y������u�^-��p��9�&{�D��J�M4œ~+6��g�����;�H6b�4g��:�R��]bw.�i�Ǧ"/�ᩊ�<y[~�˅^~	hi��D�c�,Gb!7ф��	W��茢���j�(0;hsUͻ&>�z�����~z����B����Aڗi��بt��NT��z�=�f0Ԧ����+��j� ��{�%3t�����4��{i0��T��Jd��EE]2��'��h!�-n��P$q�r���!a�C_�^�Q͢N�V�����Xi�CV�Y���!���O,A��0���OGCYX�V5�v�nc�?A�R\p�������#��rt!9���rċ�^����c��;���L�RR�6d�<3[|6o�� �հ#Q�;�������I\*�{a��Vb��%�~�
�Z�#Gb�0�D��5RJ���qY��x�T����(�H��h���>���V%�M�}"\�*U����y�l��|����Pd^�Y�:m����L�\=��7���	�;��vi�g�g�y 7��;�t��d��w�@XO������62.3!�&��;�h�kè�.N6X�5�.��+:���th�������:�?��~�ꎌ�YQAP����5�_����®��wN�*�� 1���DL�oLo�Sv���d�6�L���}�(�H5���Q�#��[�8�{��Uv����
��S؝|{>�4:�Өb��� g�� �a��oy/ҭ��K�N�Mk:M��$�_��v�Q���� ������5�}-�Of���͵�"�$-|����_�Q��<Pd��S�||��������kD]��Xf*R��9��0e*�T�J����Z1�mK���!n�߂Ml���D8 �Z�X%
�����(��I�:�$oP<��Ǘ&��:�`�x�y��鰯.;����B?����R6<sI8��ũ
!7�Q��ɘ��۲�]�Z�Za#%m2�ȍ>�u����y���ZB��u�N�8S=j�hθ��w��$py`v��r�����f��y��U��p�=B�p�y���5`�����@�_�yL�������p�wG��؆��c�!��u�r��MY�d_%�[��a<Y:�q0�\�};H���l޷�C�!�#r�
�o/��Cq5�>\+�#��Z�P`1�8���C�B]TX��̬^�V��Ye��T*����j4;��O���H��� �'?��{N�Bl�ǀg�x�1Kj.��pv�|2�����R0w]�4�f�h������/�x�����P�b%�����8)Wag���$���;��9�`�+���x��G�C�#�i����=�Z��xeS!\Ӛ	�$�(�"���ab�A4/�� ?�6���b�lS��km�b�foD�
�Gc��t_�xry�y��5��1i��ϱv�0g���lfzӏ�v�,(I�H��� ������4IZ��5㄃ �>"�St�ɀ��<�K���B��q�d9�� ��7�~|�[f�W����� u�0��ɹ���8U��ܦ
!l��>s$���b	C�L��H�l�l�I߹um�/w��~�w�[�F4���\������!�%���$QV)�I"[�!�Jף���Շ��L��T���T�`�OL�Ld��B�2uLP�m_%r���/��fQ���Bf��e�ZGR]˅c�}*�_WT9�ҿv�ߠ*��%��-�@"z#]g�������QO�a(���bvc�Sű�ï GQ�P�`�%4Q?�e[&�+<�6-��F!\$?ˏ�B��;����<�krI����,�'8Z��a`��k@Vk��!"����𸾡y�*]��cD����{�5�5�T�+��"�Qi0��ّnc=_1����,�%���l�y�y�<��ܯYqXR?����Wc������B��̢��/�0.3vp�ғݙ�g����)�T��~]�:�������ne���tdEy����`�k��a	��i�W���<e8�'SDvKG^�Î67�N�������s����(�ˎ!�^��Z_���	�j�@��.�Q'��u(�����^�ó�4��L����#ց�FDl�W�zV�F������_��w�FB�u�iG���^ġs�r.��h��0>���)�Ex�WX-t�y2ζ �"��P������i_��i�¹
�A��X�=����$L`�a����OA�PAt���.������K+
J��Z��;��[��q����	��;�
ɦs7�]�Å��|?*ܞޔ4��\@Vy7���ی|���/+ԡ������$�u��I#�f���,r��
�� h�9G>�I�iEvR��$��0G�&�BpQg��y����$�px`�i-M�� ��2i�0�����<\�ٹ�m]�1����!;�I���Ò�4�w����&BK��F�e�!�u����O����a�\c����nz�/�������+��U��o-���-+�@����΄�{�&��q$���S.U�u�9����`Y�)_�t����v�5f�E��Sc���=��ah�����\�Q��^�C����.�9�gfz�b��8�N8y�o�`o}�m�c���Z:��Sac%}Y����K�sA��Y(�3oפ���#�!�̀F|1��l% $Ƣͦ5�H���u����=v*+>�)�l<9�*�e�!-R2��N>}Q��~5:l&6R�9
�d�����J`A�7�����$�껋�F����ⱄ�!
fД��F���E8AC�\2��R/�P���\/A����G	��5��:���`�g��K�wx��k�~0�G��힛S`�afՄ
أ�}+��>zXc�s*�2��o��A(�``��,�[�d���RY�~\{Sfj/��� �>�� �d�@욒R�.��s+���S���Q��+J�ߩG��g$���je�F���2D�.S���Kup��	�����0ړr3t�4�h�����FF��t��	�jaA1^���+���=#x�gY�>�O��+���\$��@�HbO��7�����:�pa��N�(�@dx�f�@�7�|s�{�$x��4.��y����>�YM_x
W�GI� J�T��C���[�Em�,�#�4u
�:�)�������2�.Q��p��+����UR�0���#�b?ySu���AY�����5q�
������ٗ� �r6������#�2��)1����e?K��S���?�[��H	��?I��Jo`�J�=%�ϵ9�&�:3���Kc� �.ȟ���kc������\�i�����BE{���-�B�.��wsaN~�F��e�d�I�e��J.u�}���"ҟ�޶��<��8=�۔�Y^6���	�0e�^�5l�x>eZ�?R�L�c^� �]���Q�;a�S9�r�-)�s��b9�l2k�%;8U���H'�$�n�Q�Ah�����k����f��8�bT�q~v�Ok��kE�5R��;�/Dpf�/u�#�޿��|ib�t k�o�¶Kš2�t�,���N�]���^�m��D�f�a<!���)�µ'Eʙ����q�����O0�E�u\�/�"��п:�2b�Wٙ9��@Y��X�Aǻhh��Dyq��I�{'�\��eS��P����R}���+&�.��{���ȯ�n���(�
@I�L�-z��׮�t
XJΟ]X�����;G�Q'������¸������N�h$�(���k1|�S[_���Le�����j�٪�	�c	][��]Iđ��r���ps�XiE'#���x�`uQhy��(]g��l$�p�6�|��!�aw|p�7�ҭVT؞��2JϺ���ط�n�1H!�#�ɖ�\h�=��K�G���F�zq0�����!���0�����F��
/���l}�<��O5�<�[ǖ�`�d�m8^����oiSK�CL��b�W\VX�y���I�ᜪ1K�1*�c2��R�a�4J� �0+��U?�{��X\0��~��صT�}~g�1��GXZ�v��Gk���䋺�BWo��:+J*��ѦBm��AA��,���/
���Q�G�Hl�k�U���QV/���f��z�r�!0EYå=���ג�/�N��U�%M� �Z=�ؔ�-b];��6�|ëCq���2L��n2t�����*;I���X���YdacJ54U�m�'�7\�>r^'��^h���h��)�rm7sn�J� �#f�K��
�2�jA�W~M�G&G�ԍ�������>BA}��u��x /Q�A^T#V� ]�%�0��O@L�l�.��QB]L����_��-슍G@N@���pb�-�S���Qi,^nCfG�x�ߓ��1�\^љw�YAJq<«q�5��D�c�F#�N2��+k��tT\����ړ�K&*=+(U�^�D��9�����1�:����o��Se�8�	E��xp����:>��d�	�i��P���&3�!��y��k,�JA�����R���0t�u����WRD��oTaܢ㇪y�^p�,}��#@?#\!��j�Ї?mlf���P��r��0L���\Dvu�����A:�����-���[���ʅ��"�QF��狩>/.i����z�#ӶF��:'�O�Hu15gn��]lX�w�Z�	Êz��5����V~�������R�[��f�w�SSX�0z�誘)	HN.k��2r3h���a�ѝ��з��u�g��>�'�JtfR$Aي��u�����P�u	HK�_h�-��&˖&�\M!�F|GРG����s�V�	�����#��e}6� �D� G�1�;"|�\PCI�St�������l����>�|[/C�]pw���w϶F	�'�Rfv���X��G���Z�H����_�[��W���c�IPȰgWt�)"i��R[��T/#�H���9lVst�T�S���N��Da�UL�HG�[eUoGY�?��P�m�6�[�j�P�@�����z�Z���Hm�O-��	����B�f�:M�@��Q~�΁��{�~0^�G6ơ���-�iP�� ����
,"lpzN������iGK�]Ei9T��@c`�z~K'6����x\����5r���_I�OF|�1v�^wtH�le)~�`��vQ̵`�(�	KL�˲���"R�}�P�����Č
8*��[�<�́^��6t\�?���NKv�6/q�ۅ�-�mXw�C p�vL>��P$2-��~��v�2}�����R *k�ӢD�?��O�A�>�(��UC��g�F>��<Ĩ��o�a�����r�o8�a[�>Q����K ���/�_�eQ����T{Qc�;���K�>�MU_��ac`2��Ӱt6C�;�c�j\nNE��c�3����Q8�,�3����3��J	Z\0��$?�aa�W
���UCI����}��~�nQ������6�ށhY\>7�
;�m�����7�
���w�s��F[�!�SQ��8�ʞN�>��i�X
U�Cj9�84o̤p)�����H���NFH[�Gbe�l�5����u`[����*�wi�W�[�u����gr�s��a��ո{��v|���W-�&��c:��]"���^a�kG|�z��n���GjC��������=��E�t�@���W�߉	����B��yX���?�"�1�mW4Iѩ�֟ú�)I�!�
��d�R�,�MP\� (���)O��k)*��JZ����b�I�	N׉��@h�[z(}.�E�#���Z�������j��j;��z5Ci�o�5���fl�� ��Үw[��3�>i��ƈԭ��2��*�9�G�6�Sa�4�繬{զ/#1j*wU�T����&�^��B�b��Ŵ+3|��X�X���)Ƃ�Qg]2'�H�h����y��9����P����9�D'��w$Խ��d���@b���F�ٞW0��.Y���*\��Z���pƃ���3�O���zZ}S=�np2 �N`[��_���h�1�����G��EA��K�����~�w��0��,`����4B���Uo�1�P�,ǜ|F���o؎�8L&Q;� �p��Щ�UgAw���ϔIt��6�A��h}~L��T�dQ8���mEE���O�Ar<�2(5���  Tʭ�3VK���`K�L;I>��س�Sj*�0�u���+�xG����K��oT�����5�=�]o&��1˽��������)[}�|l;�ې9Mh�H"�i��)HH0Y8�<3�f,�نp�ThGw��l4�R&W�:��^�IVSi�6V�\㧞�6[��<ls�v6 m�ܚ��n���R�J��T�e���y�mrh��
G�(��`G)=�*� �R�'�O��^��i���G�H�7�f��	���b��$p��!Z#�)��pK�-�>�Ո�`6�� .aTu���v��2���Z��G�F��u�L8PY�{�2Z�&A����?u���P�ʻ�Gl�UCG��	J_�']���,��7;��L���1@�W�B�n.1��Z��s����؎���e%��s[�N�Y�JJ㥍g'_67�-ٰ5�)<������=�n�C�B��c�]-q�5�%^���iy[2<�2�F�MP�`�A����F�/9n=�w�	�ؽJ��H濊z��\r��1�;z���6|뵿w��h'W�z�p�a�!o��R�q@�p���ջ��׳�:׷3���2�}0)rx����g�i�!ƘS�{Z�m^]	�1��k_�L��"��z�
�ґ��\����\����В顣ӛ�VC�GkW���ͧI|���g��!lPtf#ȏrk�!!�L�NV��dˋmh��T���Y�����X�4u��PP�Yo���[n�ё
'P�FO�tOx8��&�I϶���ttY��#6Hk���ۻt��8�o޲����8$��n��U�W;�8�Į�J�K��k�Z��j�&�_���4HG�c����q�	���K8��u4�*o���3�Τu��P��qQ�1��I�T�u��������94˿���V?IUu�Нʦ�|�i��T͋��fL�4�Ɔ���Ӻ^���s�o{��%�i�,��Y�H�(���}RxT�m[����w�)�'�k�LXu�N_���i��fK����L����ׂxA���<�N��(���N�n�uzx���VՀc��x�mA����x�,�T��c3�~���V���a���
