��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s<�i��N-X�4Cx�û�M��TH??�[~Az�?�7���?
�q�޲H�=u�^��� s�$Z��J*�wQ/Q�,��[�h�s�B�kUq�3MQ�����>�j�M�,�,���:d�3�q�|�����5��Shx���gy��57�ǁ����)���}�����+�@	(�XT�M�)�j$������ɧ����=�H�e����ٜ�'��>�u!J���|������h�?׎�r�01�C�eO��^���E4��I��g�ҀQT�y݁��Pl��\񊠉%�U�T���d�э��(&��|8C��##�N/U��"�;����c��V��i&�j�0��r䄰g4�s:6��g�+�uv���R�7m�2G�1*�a�u767>v��4TZ��s1�T(˜�O�\^]7�p�JK���U3�$��Nb;��/��mN:��f=���qFẑ�M��}�w��	eO��߅���N4��
1�q�����I2�&Im=�Ulɿ��fq���m.}�V��I�A�nTٻ}�ղ�,&�r��}TMWj�~�,�S\��N�-�<>��'��������]#�.���-;�d�Sʷ�Ō�#Dk�����s� ����>��ޕ.���+���ߚ���<�#��Wd��p��1;BC�BS	53�i�d���^�Ԣ����DV+�o�Fd����YF2	� ��`�����+��
d������p}8�U����]�헿�� j\$�)ዎ�I�94�z��+�k�65i�R�
3��t<�#�UKFӍ�1)NKh��Y��jP���+�[��7S�N"��}'���)4�u��k���⠾A���Ps�7WG<7p�{g�������hҽ�G )���c�[�-�Q{�٫xq�#^> ��������C���in�=�A�XHj��xW���]dN�`�=���u� �K���ý 4��i�(��6��H���k2�V�멖�#,�Ҽk���~Y]��3�&9eO�c��U�#UgE���(n�|���8P��y��6� $��=�{�>��?�+�<JS�K{� ��A����VK:����g�i�{R^��SC_4�!�ޅs��Rm��Y��VhG���34b`�\$��No�/dȑO7b<<���*}����{�¾E��;���s<�|7s�U'���p��9i�I�#=�/ k	]��4�v��q���׀C�c�|o*�s�ƅ�fq���c��յ�q�+�0�
���	�i����2e�*\�JD0G<߮���h4�T����Ԍ]r�(�[�����T�e (x�C+�����߆{�?b׺J��ak㩜7vU�;TXwg�,�a���hp:w��o�1�K��2��
Tx�T5 X�%:����q�Zo�2|>`t�������eԭ���!��($�}��Q��S��ʷ�;�dT�b����X��YƇ�<9�1�s���	�=����T����"��Bc������g��MZ�<�j��޾h��$Ր��v:��� ᩑVD�y����{rD�k`���R�"h6�\��U���j�w	y�ʗH!p��?ss���� ={'Ji�R{u��~_��?���x�Z	费s�j!��8?;�P�Ų �_n�YHfv���\�FN'v܁���`P���@�kb��F-C���M�����J�|�x������ޞi�l��d�R��'tR��qx���8��i������W�w�V8i�{��̥|�q 8UZ8����Ͱ.=�ܚw_̲S&����u����6����絪�4�w�W�z 
�	�c*:`Z7y���M�f�r�W�a+M<w��ލ��O��|�ܻ�V������u/��Q%>��i] �ߐ��>��[?��i�#jbUwÕ}��Z}���X�s�y��:2{��2�dV���7����2)��l��� +�ѵ�����pn�p�SW|����$��M��v��ƐE2�+�����!�J�����;َ3�P���m���M��j-k����M��ב�j+f@��n���Ҹ߁���J|�X��FJ��a��#+.a'���=�4ր;Y�wD�Z=��VU���MG��a����nT��p�C��*9������K��[�w/xt�nZ�I��|�Ge���`�_'G�[R����ﷳk��T�D�'���*Y�k|aL���񅘊�5�Y�7�oI[5�	n4ʦ��T��V/j�'"�D��<�@�K���2�l���҇�؍�U���~��B��p�������ݿ�%g޽�\����N�9t 9�U�<��f;�rN��<v�%L`�:�d�hõ[�1�!L���@�W���3�SmG��8޳�<7CV#�u���B�����M��?%�Q��ܽE[8�C��TN��I@RɆ����h2��6���Vl�/J�95 Vl	S&���Nn��7������CZ���J��9�ϛМ�P�77��5�]D�o9�©���b�(+Z�wޱ��r�8XM�/PK�՛H�ScU������9�s]�(��4��������
�X\�'.��\�\���;~�ֹ���i�e�pv��wM'P���a�=��µ��^����LW0����mC�t��]-bQ��z�6o7����I�T2	W97L��a��p!���謀��D |h��Grqm�� |������5b>�N9�xe�N`wf T3d���D�;�C��m�� SwWĺW�ԡ���Rº$<d�,gcO��������0d2brR&�����G�%��_6���T����?VD^�/9J$��c�9�S�C*B�5�~���lp�`���t�l������	�\����w���f/�-�lLɎ=��
�4��	�B	��[�(%"5y�AWSF�Dk
u62�A�܎��a\B�t\��f\5�0�!�m��?r/L���c�D�?��6���T����(�4Z�������V�GQg�Y�* ����)�g�D�(���]ϖ��M��6�z~��Y7j�"OQ��l%���Ql
���i����-�q��tD��&��a؞�&���T�P����z����|������i�y&Y�k�̽δ��X-��J�d�>�qBUcl�6g��]�`Du�(���ܹ7�R���;�o���QO��<���Q޿D��Z*���U�7�tk
��+8�,N�M&�������~X�Y���}��Po
h�H*k�������~�*4�[�~:�Ȭt�����"����������3,h�-���=^'��d禕?.A�V`z[�oW9��=�<�����V(R�G�@|Ġ���U�ᱞ���~&g%��@\�����4gפ;~��qV�z)�=��1�;c�4��>��ۑ�d���D�l!�6؜[[�������]1�,-	�����~5�$��=�v��Y���h�[~�H!dgk����AG�t?_��n��?pmE�|	��tԏ����Ƕ�TC���c�����K6o-v?Zm�3{�������4�*J$aI�a
��=��&g� Ko�A��.�ܘ�E$ʤ(������������F�J�J���S%6�\(7 ��W��,�F)�R?�'�+��
�})ru�VhCԋ��W���R=a>�߬�q�¶wJ��D\��k��_�ڗK<��_��@�v�����ܲ �@�]5\^	Jp�#ɤ���_妺_A���`���X�s��Z�������<��'R�lf����=��',�����k|� 'j�@fy���e&�6	��%�R֍>* B��l&�q�`��Zc�}<���0��
�����(��!� o�3-��OF�� ��Ac��D!ͻ�X�zQ�u��t�l���h�W��`q���!3�Ekokh����#��ۻ�Q�u�-E,R��H�n�®9�m�#�ً�AZ��9+���iQ<Jl�^���0�ϓ^7��� �F*���(H��u��H�k�t�p�˩9�:�!U�T�E��E����{�x��n�cd��y��������*�D���I��Ry�q)��2g���lKVZxK����
|g���G1.�k�O����=0�Մ��� ���1SC�cE���G7TLޖ����h�����y�sS���5����	Tn���n�>Ito�$�H�^*9��������0��;Y��g�y��l$��2�0w)~m�8��T.?6�)�W�I\�A4UL%BD-�9��-��>Zg����@��ټ�s��%�ߖ
��M>�4��
4��zǘ���\����m��D�ʉ>�����x�٪L@h�ǽ�7kD=���?��u��0uL'|�{>F���Y˟����W�Ń�Ȭn�42�Y{��<�9t��<�"t\���F�4a'�O^k�1�}
�P���8���,�����=����%��qQ�n�N���g?��\ aF��Ա����M����O��K%\`c��<!%��WE��Y6�:_��,A�uo 1F37�t6���D�c�V��� #�I���.���^8�.>�׉ڇ=�k@0�p�#D�f���ٖ͡6�$6�0�*�72ŧ�l����<F�l1E��N��$�@c��*#k3�L�xB�#c�=�;��C�l�� Zc����â�9��󏱾���z��[���,D�Y�K�#r��;L����UkL��P�Y���:mc~�~� Qcˬ�������uXa/�k%^w�4x� &J�Ҫ}�2�krOV��ܣ���^:��5� e����5Y�F��s@�g�y��
K�R����f��R�B�{ ��%P�s@�B���t� �*tu��N�5�6��6i��$��tD��Z����v�J�����TL-�ύ�n�#:S\�9�����������;'ә��7�-)"���^-�RR�㹁���aA.d _N�$������7�_6��iُ�y�T��`Xn!���K��+e���]�Q�H��/��(��D��%(���ΟO�B�J�������o��V��p�Y3�{�KlѾ8����PV�pݭ��X�*���Z��}���]0�f�})g	�'�BGD<s�?O��nW�	ۗ�����=DK��=wvE�|�7�&צ�(? #UW�1ԺI=`�,����V�S%�	�GM=�GX�ro��a���j�������+M��
��1�q�J�ȂpQB�J�yˏ�����+Q"��\ƽ��$�Y'�D�����L��)�P��_[�(GG@�W
���cU	��s�"V4K�u�}T�/@yΠ�v�U��%E�v+%v1�5j�g�(�S�tz����Qfl�*��G�P�I�y�w����|q��t_e0�d�Yw����ނ��8��e1�͒��W�M���0d�xÃ�)D���� ���Zl^Bw�*6⪦��X�(.1l�Ȝ�O(�N7��Y�E&�:^��E��9����������S��������;�o;���)��8��|��v�h�݈:�ϰ��%�rtu��=EȈH�T#�bk�����e�#K���Ѩa���	�&�"��c����o���gq���	��p�Q9���Ln�,E�.5T��ܖs�c���N��g��}(��l�7Ex��bЪN�r�چ}��
'�L�ܔ��ල8�����:V�[=){*~c��R?�-l^�Wa@m������;��3�����>�zq�Ykͱ̱)�i'v��!Ί�W���;>��ϵy]V~���r���!�_]�j�Q��x*�O�>�ܤ�V�T�&9W�q�i�4���������W�P����o��&E��8yK$8�[�g�SHN`�'a��j[�Q��u��$/��|��B��ġ������V�?����O�R_v����ě?�o��]
6��!� ����O(��Xv��3‛������?�#&���7�Ɠ�&�Xg���h�Ͼ%'wXF�j��nc���!���&�8�]ކ2.4U����Z��!dh�HK��B�N��5欫�^$F:�O�%�`]{ЦE�kڽ:5��o�w��(�6�p�-�/�m�/��RQ�6D��Š}d*D�j�E$�R>�A�|��5��k���b���:xp�o"݃"i>/O3��ꈨ$ͪ�{N�c�>Mx�$!�S/$�����m�oL���ك�̓2���.+�g�y<��E�'Ut�K�@�����U�b���h�*�O�pk�]����wз!Qy��bb�e
���l�`�YW��&���ǳ�+s@j�4�l����[�L�9X�s�-�-n�w'M�|�l�9v��'��~}N�M&��<�,G��u�{$��]v����#ɻ�m^=��7���k�ʊ�z6
VH�V�֦�8�l3���DN��I�������~��_D����c�6��(�r�{�h������^+
-�O�ye��]L L_9��Њ�K.��g���͢�V��p�������@��)(��ENO5�t=���`�qʠ�!��M�ڻ�G�P5ȡ�Y ��3���pr��B/���Ga2�y�
}B�nE-�[��_W b8�Id�c��aS^Fߺ�����Ԧ��WK�g�X���w��ܼ�	�A���kZ��߯��r
���ט1�'�dr���FJP�":Q���N�X���P0O+@��.9����*�5k(����r� ��O �D�y����]󰯦�PS�w�ru��)9wN�b^x�Z(n� �}qL�gT)�f--�/������+p1�Ȕ.��1K7����6��*����S��j�y��ý���7�w$Ħ���X��ER��w��N|Z-�HgN��Z#���P���t.�+���g;��Z�#'��.[j�lĩa71G��\���6��˽��@�x��(&�+�+G��IZ�n,�ń���� ����ҌQ���5�iWY	k�[@��3��쩾{�%���?�
�`"��;4���~|;z��,ȡbX���b��`l���K�z��]o�z�9��%8IB/����@�O��s�']�fe/��r|��W���� ߍ���X�G���_Y�n�^7x%H�J1��|��!�#8"��o;Pb~>lc\�O � :#��|ֹG�HѨ�)���G�F4�.15�_�µ����$�&�e�ּ< ��4�.�_\����6�%��h8��&��q�|`��6�X3��K[�Y�a��>K&�V��M@ł}�~F:T�K�@�ޑ�vbEڭ�WJCBë�� [�Db�:W1�l�a)��:��D&�)����s�>[�
ZЭ�(ua�{���/1�'l�;"O�����붌{,-g��[;��Q��۰��}���H;�|y��z[��f�`�Vl��}G�"/?ރƻ���ɎOb��?)���5�n\�:5|iNP1jFc�W>�.��;��6j�m���^?�������W+I�B+�3v���؞7^���QB
z�U�FG�~�-��~d��.���9٠�%q:V&�$	�0��H��b�_*������X�����)Y��"ZH�s����l�����$7W ����Xl��!^�_l��k/&t�	�6�1 ���} �W1���M���B�ó����$)��y@_�{B|��d�m�V{(����l8H�~����@`�{��s�ڶ����n��.Ʈ�F�+�)u#䦄��iJ����`�p��F6�i�ɘhl���"y�k��K��}�_֧�&�T�li��O���LU���2��2HW3�&y�G'B�i��g��Ũ~P���Ƃ���gFT��b�*�褤�j5�c��;�� w(C��Ew�ɘ�w��	5#����g���3�uX�ʛ؏��PI'�1�z*�â��*�����%
:�˝�Er�F&ǭIq��R2Fئ~	�`�ᐾ}O؞g�xx��ˌۋb����X�v�Zz��!�K�T�t(����z�|1G~������`9'��2줵��Vg��x|C
�jf�\�(}�Z�l������1X&}+��پ�����h��!le;UN'�{���i9������&=����Sz���!/����+O����,B	?��:W�|����_�Qǣ�UtD}a��R3�B�֐�|�;��/hj<B�Ϧ�	�.��E�@����6��U�#�K��1�~։/3
���窽J*��&�O���E`��_���S��@����z|=��\P�[��)��{�n����b�Dӛ�@�����em�����t�e�������e�$r�9,Pxf�6t�_��@��*�:��<}���b X/_$�m>NhP� ��q�Bq�݀U[t�;���8�r�DB���pQ h��w�?"��ڄRPX3�s|i�[�P(�"Sp�wr�v�.�
l���J��S��F����[k�mѠ�TqF����`D&ϫ!!��+� ��6��PV~/;�%R�� ��Ǭ�F���hD}K��<tP�r8��Q��g����� `4�����T�e�cg&��lW,π2k�^�o�D;��B�P�\\������d�gN��ۏ<Y'][�Xtfn�u��30��F�桃��0*�|��5�Z������F�_G��Y�%���k�=�		���ׯzZPV-�F3F��{��`�p�R�g����a�%�_�F��1Q
	���y���������ULc��iF�ip��P�V��@s��vS�ʹQ��D�O�>��Z�	�/����F_�7T�����=E$���S(��6}�̞{f�N�����U��;)����fts�4%ʀ[�Cl�D���A=>LAc�1��}{�OmA�h��8k�|��֮ވ��7��Y�3S��4�A�d���g�H
!.�t�HTV�0lY�_��C���,;���~�F`����e�&>���-0�U��O��~���zpxXT�$��U:�
ي��\��&�A��z�J��\�%dPo�!8�ةܝ_����Ȩ�r�n�wã�"��B�{'�ă��fN
��������'	*t+��Q\x�ʘ߭`�����s��e����	k�tmW���z�[��5�"��	R����m*-˩�K/���˪��md�,�Xt4Z�0~tȴ?q9��)�~�̓��N��Hm1��]�2�n��D���Q`���&���ݝfw�ge+��cʥ����}��8�j��:���)�#i�tW�K���H_QH��h2)S��L�t�_L]��O�NQ����a�#���J����������\^dlp:��p�֊|���^�F�>yI��e���o�)�u��ydr׃�(�<_Gu����}����o������mLK���<��������������y�V�e�4X<��G�Q�%t��H�<���Rb���3J�<?$W�GS��k��LT��|�lB*(�����j��ĸ��I9�h��!|��s�3���z��������B�ej�S�W�KG��;�-�Eq�'��D�	�}��-?�.�&)<���|eꇯ�Y��Fr��g�`�ٸx�\J��
