��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��I��i}6�_��Rf3&q%0��-��/3B|��P��Ɏ0wk�N�Fy�p����u ������cS���ԸV�z;4kƮ˴V�:���]8j
�,�YğPѾ!����M�E��������eg�RV���_w��f,i4	�����0p�Lܧ%}��떁-C�F(��~�ޙ�����~�F��-H�¨�vd����n(����v����6��/̇���ҮƐ�wt�)w�K���;�K��JP����
���~̔�b ����h�]�kGtub���&���h��5{��n����CەQ����� EM�T�����H�?B�/^�Ӗ�'N�
�K���#�.9�C�x��\f�~,�)F��|)m�u�_F�X�gÃ
��"7y��-V��c�o��o����w2Zi���S[N.?a`�[7q� ���N�Z�G��X�u��	���
���mx?a��x�O��j 6$/�v_�{VaL; �i�WH�CGl�2�R�5{�U��������y��Z�]�k~�����R7� �Nv��R�p��3
��U�8��(��'�V�U�#�B~-(m�D���K-�x�|R����C7e���U�@Q9oީ���xHF޻~cA����(�xl��ش>�}e�r'o6��|�Ŕ�٧���AI9>:�EU<�HV������D86��x=��ڮө���:yD��zߧ�!�1�
>�I�w�l���C��9m������2^����DϚ�����	�Z��ꂄE-8C+��� y �^�OY����Q��YU��dh*���$���[K���u��љ��^`kip�J�6͝���Tf���yzN<�1�.I��¤U͆�#_"�+4����DL����h�.ow	�tV�N~g��i6l@�#�~�nW��Y^*�
O����`V�L�1~��ڨއW�ѱfPEE�7A�7��O�K<��@*��a�����ˬ���e��b3Q�����7+�0M��4�
�ƶ=�Uۍ��!o�r.���Uxҳ�v�O�v�;�AD|�q4E�á��+E�^AsRhhd�����z՟��[�ɼT�*�*�ҫ��ь���i�Z�[��?��W�2�w�S/�w-- %Y�*�dq�!�|ث�Xh�`e�4��t����F��2D�D{To�È��uS��&�T�+���3�T+��������7�O���Y���Q�'���`%��P�&�u�;��+ĭPp�3�dP�������'iR�bgh7�����`^w}{��P@�T��u��"驊����I08mHn���1��I6̯��DO�a��BN����2"y�·Phx q~��8���dp���l/+
6����{���E"/�i���aT�$<y��w/����k����"~��/n���5+����Z�*b�!%�c�������F�z*�g#c<OE���r�
afI�J2�#b1�W�d~�5��5�^������U�.����ζғk�����	�I����٠�-�0'y	#�-K�/�Z�1�<1%hT�v,J��j:i�0�x���W3m.QN���֙��Q���w�� !�H%��ڧ��� �ʹ��4#�� �mRr�R��5*x'��سrBqs#gpL(��/M�O��wS콽���V�"��?Z����������<C��Q����Y�9���t��]޽.�%:�7Y�]ܧ2O�o�TM�ئ�Z�"$���7��2	K�&�j�q�c��d�@�::�$���a�{h���%��ݟB��^Sx��Y���s��+�m>�8�����D���ϑ����O ¬�B;�&�>[������c-4'R���RH_w��7����5diQ!�D2�������̷�m7�A	Ƕf|��q�Hl�
v=�'��1E��1w[ϟ�X�ȖѢ�6��� �6mDk�$1�������H$ ��GՎp�k���W�bzoً���f۟0o�lS�c�
���,���u��� b���9���z�� r
%Ĭ��sk�L�5?���l���r8!��;� /#3�ng+��}zx��$SIBn���x �`�o�``�����Y�o�h���Y�������{����h���i+��6g\uSP'��%N�pA��ei�����_Bi�1BՍ�I�*��7�pҕ���44&u;��9�|��b��6V�T���9�6�]^��0� �=��;%Hi��W<j԰ƍP�Ua����]7�|$��)�#��NC4%��_f�	��h���K�s]}U�������$-jH*�����t�P�?�	���$ݾݿh�x�Y��rj�_�T������hG��f�7f;%���fbݾ��Zm$z����Ă�!-�.���ڡt( U�ڲE(~�~�-�L���E%2�K!ȗ�ƨ�K�t��� .V��i���*ؖ	�	nWױ֥Js��3�Ŕ�(i�'�O ^ַ���H�̦��<I�)��}sh=��x�X�	���!����U�0���w3���~��+5H�
�5&�zO�Z��G���G�������q$��c��ŞT��>	�e.���y������w�������*��A����K3�x 6�sT��e�Ӭ��N�87��ޒ���%ff��:�}\IW�f�z�5�^է����,�~Ve�+B��j�cH�|��	�ÉJ��3�c�n�7MDUe�to��بǟV�� ҽ�4��v_�L�q#�;��p�\G�;�ʬ������Ia��D����׀��bk6����XY�U�����Y�Y��A�H7c��g$ѯ��.q�8���r���#�D�C1��XOS���|�2��v��UH��L��ɓ�~k��ҿ��vbo���j�+&���ʈh��B��p���E�{�V�N��}���-��S&�Pd\��[�\�8�+Z�6?�kd�oB�?n.It���� �-@��{��6���3Y� l{�U����B�DX���wnޟ�wU��O�l���qH��rʾyA�0��.�|�b�Cǉ��%<���sk�ž�WI�D�i$s6~1�e����8������澟�u��3��̞�x�L��*�B�RC�H���#V��i~F�M���Ԙ�E�)2�x�47��"YB�ȉ�j<֣�Ð�
�K�V?�׫�Wv��ih����PG�6Z�������O��1pl}� �=��(`URf���p#
�f�Ѐ�����j����-鄝�1�L��7l*��U��+�4�3���_�1'�ĳ�����Nz?�" "����н(���tV@+Ǎp?�����s��r��ٔ9d�}{��ĸy�"�(��ǁ�a��D��p<l��1q}JW�4���qH+�nɣ�Q�O�G)�YT��j@}�����֥���ן+@�	�q ��V�ID��V" �cl�A��e</��(�j�0H�*Q�7dD�'�S��5e�}}��ʵ �y�bzߐ�D�K�W���-��dŋ�Q���-:��OED6��?@�Zǜ�E�2h����#ӌc.'����P��Wf�8*�_}��h����	�8n��\\��uR�d�X�2z�v�=�>]\���)&�0Q�
&9G^N�Dr�Bn�\��g��C:㌰��)Q�]��pF0�I�2��U�����0����&� �\|c6��@��:D�����f���г���t�C�&�a������!�#���!��on��;��#�}��'"�T����S�J*�սqflA1El8��O��[��V�ƺ)aX�Te^�����l']�$g�uWPn��P����+e}ߛ�
x��x=Qֆ^�r"�g7.lCZ���E�E�1.��P
ewu���mw��2�ݺ�^,�6��e�.t��88���mQ[��?��K&�=�ޮ`��1�$�2�C���@��HAߒI�X�S@�;�=%G�:?H�\��P�\m�ۣ�#��a�<.���׾�5_7t�˵�4N$.�[�蠺9p�Y���cw��#.�v?�X��Bm6�����d�����4��ۥ,$�I��������w�㑎���vl��N�keI�79	��~M�Y�e�F���{�ʂy6_@�[��/'Y�anPn��	ix��ʖ�0�����>��R�*���鲅���}[c@r%�v����Z�.�s(�jN��_ýi�j�L�`�A�n��e��No�y�[ټh20���BH2��<�l�+r�gE���Ī�F�]��[�qק����^�	�>�JW��=�Q�i������7f�pJws��ᷭ�v,���sj���R�����vlB�9!S(�!�]4�P��3o�urc�����q"����`����g�-y��w,�W�J�)�����#'�ׂC_���[F-Ӷ���D��TY
�Ye��d�$�����m�+�Ի����8j����0��=y⾈8��d��C�8�Hĭ��tE���#�XtM
�@�� �B�%�޲���,���Jfޗ�&��'} �P��7�ZT� ��d�����`���XuҜ�T��#>m��m��@p_�՛9��"���df�����\Х��b������y��B����x?�'����cI�P�3yho�������S��8�i��b��K�uNx柬]��Jd���.���q��v�B�n�=򨗲���'�س�Et�f��B�jn5�9C`\����>�0��ʻ��\�W���o�*=	��|A������'Q�J{E��t��a䟑	b�s�@u�W7�/i2�����Ǖ�w�Χ�r��/`�콟Ld��rw���G����D�_��	/%O�U��;�١��\�
���,���"� �Th7S��.���Z�*�/m��#΀ m.ΨŻ'��3�����(��7�7��P�4��a44S���7��$^}����=�!��L����dc�1Ac���*�R���?j�ook`0�WÿO��:&�l&�����'	��@ǟ��V
���r�Կ�_�/R�WK�y�F���{�_lp{��i`��14S~�a�����r�v��pF��8ɧN��E���ki[�]�5M'��+�跙� ~0zW�8jݪX+3b�oS��Ri9��ꨏ��T	t������#�$[��Z��jm��c�z�1B����{3�p<���x����������[i���A�B�8s�s���فA���w����y�q��������]���6��������T�;���j�qn~�� ga�ȀNT�~Ջ+��r���専�����]�\i��
u���^��6����CK��#�Y�GԊ1;�pTU�B2+9�qJ\7��	u�
W��!r]"o��w�tޅ9@x]F-4K�j	���#���d�o�l|{=`�P\q���	t'�[�qׯؤ��SrB(J�P詴�����t��6��w��3�����L7ǈ[P���5��'A�qp5��'�]���ui:�39��������t�!�}���5:�����?}�i1����W��ѴK%)�~�f�e[�Qr_q�m@꛽(?� �P�T-�s��0T'G���Dn�M<�&㰟N>���qoV$����/�pWV�t�����?�XU�@�5�0��Q�>�c�?&�FM(|���9҆[�pB{/Ϛ�e|u���N�@�S��Dڶ
���*�(��,�.weS���E�A�D�}�����
��B��zFN�q�K	bE�����a#�i�����Q��9_ٟ�I��jཞ޵��ա3�	�?�h��s^���j�(Bf�M�Xު�S���'�jxF慤0�p�_�K�D�cx��,h��g�#��8�4v]�|V�Gf^�˒#�s@��J���t��F{� �]��Z�
��UVrn�_�Z���d%���quH�m(������7��K�3�?�Ï��Q��W_�G%�A�J�}�*,���,'����rK��&ã�]���l���^+#Yz���-u�FJb�(8�����d(����R�](c15ܾ����Uu�T&���B�cD�'6
<����@����V @�	@+�-��ё��x{�za2o�.��lm��L�z�{�=9U>����~�Ҕ�A���?��2��:!���>�G����_�J�{i��aoCM<��k �|��6��e_<]�G�;:d�ǯ�._Hv��}���qG���]�JH��b���i����5���o�:��F�s��N�j��5���WGw 5Y��,�<�Ā�?L9�	��j�}�m9�U�SS[[�]Ǜ�]A�Yw��|� �Nz��'ӡ� �l"�}+1�t�:�U��k^�V!��?�C��[�������y�ո�}�E�̭�<ojI-*T<�P�i
/�~�E�rBu
�S�<ο��^s��CA��	͈��e���..*M#�ֳ�y���0�:�D�C��@S�g���[S\�M�p)�l�&3ϝՓ�+�"��ێ��#!6m�3�ճ�����X����m�4^O�CL����s.��̾d��M��0�G��Y볲K(�-D�Y�ѿkLL���N�g��[���Xy���7�r�'z֒5Z��3�x;�s�k����4�GO��uiv����T5����k�R���O�HQ8	,�	��,��74d�'ha�/9�i#����Zř-T#P�����|� '�B�Ǹ��C�aA:���QںI����&�/5��}�R�.���tq��>�Y�"
H��s�x5-����g/H��E��� ������Ȥ�ڶ�2ϙ�k�˾�!��{-f��L5�L����:�U_�y��_��c�m'+���r錝�\8��xU�*p$1��?���E.��CE�8d���D+��#;2�f�X�ލ����8���o��EY�, � ��O��(#���;�	���� @�@�;���Yk�"��)^�Z�
��d2��.�ܡ�u����3�yߨv��F~SR�@-�g��G��<�$��w�H}��z����.��e`H�.a&eѕ3Q+��Pdh�=KR_�|tXٟI�t�X�

-D-�G�L����ٗ>�pU���9t���KE���i��gۺ�
�5*�e����r�G��(�s9�_�<1�-�i��A[ �/$���P
 ��T��	�SA{w�n	BL����.(| �Aρ}"��onũ�t-�(���T���X�J:z2���z��J��� ��,)�~�>��2S���d��R�%��ƪ ������=#��m�~�x�9�����%�Ȯ��e	3u�d���>�+ق�>��{���EٗC����g�Ԉv�0���`=wR� ~��t=I|	|�*��/`�͡Sp�0�����%x�2xh�J��FWt��������ͷ pG��$��/��~hi�cSq��7������c�~�G��(R&��A�ME]����r�D��6[��&f���Ϫana�S�
b�d���#����B�:N�?��%��I�Cg���>����c0��o,m����P.f�u1z�}�Lz�@�c���h���w�~��������h�$_gŴ��YD1��
b��1���I�Tx�eC����t������]݌�$��Ϥź0� �I�v�#J;6�pBM�G8���0.�D%mkMc�1���z�)��Ѭkq�ҹGZ�HW��:��Uzm�B��Q���þ��-�l���mAFd���{q�o�Ky�_<W�Y|�d��%3���(n\jy�U�u0iv�����$뿝��ߡ�Yü"� ҄U|.��� ���ȱ��͕� S�����R(�dK���P� �Xs��Ф2
jb����*������V��-B��>�c �u�B�Us��IWR����k�T6���c�G�$�2��+�9��Q�(�#4>�b�/)���i�Y'���@��h���%88��ĵ��ߌ�p1��M�i�;�@]��BrB����#��f�X�w�Ͳ���M0v®}��2�Tx���`0�Q��d�(�,��W/ �&-������m�.z�l��c�F���n�+[T.�j�A����OO�s�v*["\8�4�`�������M�-C0M��u��șd�N�r��<7fZL9����Q>��Q��
�X4�5�{��L����O�����	��4MDg���
d��Bǔ�C9r���-������H�W���P�b�����]�+=hxTAq�`���2"O��&���M����Ug�c�g("2٧��}��0ƒdTM�:H<��{D����=�������aWS4��͊��15#9��l�֞h�(�Tj�,���^��UZ5��o����C<-�Z�HS�=�!=D���Kf�/է��ء��kui�F#�>t�D�F�u���������VX�.���$DR��f?�ߪ�j�VdAo�3�%��y�Vq�W}��7�����%�2`����gܷ��cUc"74�[I�� L1IJ�L��?
����t<��t�� �q�a�j�v�d��3��>:7����૴�x���K&�1���MM~ݿ;������ҧ$������J/�jY|1��a�j��_���\BH,�Y�!�.��K�뵨񅖭3�\�+�]*���oK�:�M�sjZ�GH5@�k�Բ�Ԃ������,kc}pm�z�+�!b�#��q�(�{�m�2���k�N���+�7m|g%!ʃ��z�6Z"Ϩ#��C�[](��}������+1!�çl���ו�="Z���EO��8a���D�I�� "��|��6"͢��"!�|�6����rf�&ꝊQ!����͚D{4����8Or����2�'#�؉d��T����MG��[��?NR}�t��Y�R�����������6�n3+P�fܑ|.�T���������z�K~{f��j�MJ���/Q:��V����X�-W�#r��6��Um�n����v�#��*��ni�)jq��?2~�J^j��Y��m[�B�E���Hk�."}�'6ڍU��ss�,Q���L!�B칑F��-$3�TJ�j:d�u�ˆ����i������>�ĭ��۟rGΝ�Lf1W�Fh߉���
1��c�?t�/�Iϖ��'������>�vO�K���2���٩������c��!w�a�7h���	��WAb����世���1zk9�e|R�<l	s�M���cP{�� f?8v�7i4֕�z��X%�!�\nI~�uqȯI�y2+-��ٙyKD(����ݽ�Ε�'0S��u�G������`��NB���?�K�.sLV�M�z�;�7;D@��Sg�^�Jb(�~N���ēw7�n>ͤ�'x;�՛bF,�~�k���_��e�p�*o6��0�$�N��oxef�Mt^��.s��:�L�j/��e]s8e;"`o�0�$c��ԯbu��L����G�����Ӧ��}�����]�T����f���v�+��md��
�.6���e�}�WS�V�]J�@�_ s�"c/�m0T��4�./
����B�4����F$�"�C|!&d�^/��[P��`��_�������*܋ۗ����<#(O��Q��l��+g]�&�C�Y����K�%�|A�d�3����a����Lڎ�a5����ޘ�!����FzU��^$�XZ��1D�P�B�d���%��H����xAAʙ5�*�����[��1�*~�f,�N�5Guʖm����E��O[ c��b��c�=���Tyc�.��]����X������;��$�<6q�� �c���)�*k�|�o���\N�k5Ov��� I�v-�cܯ�tc{$��9��������K{��#y�.�.F,������k9��:�;D~��"��z<mbb�9q�I��ێ�B��Xؔ�>uO�="�Z�����EDq��<p×]���
3F2�9F��f����"y���Oqb��}VX=ΜIʯ�@�E��E��j�����gex��Ī�F�PO��*�)~��{�Z8@�2�(�7��s�1�eX���|6��zF��4�������g�ݷT�D��f�����B*�L�E�٩�Z�u�Y��F��*��R�H��d)���h�f���W��x:_�Y��o�4^\�A�:g�/H��6�8���4٠�8X_����ּ;q��y���<����	yXS:�k��[�\G���ik��ɜ'M@�6��׾i���J�iɓ:_с� ��UC�%����*oa��q_o|O-�⺘��b�8(`KR��vh>UJ�/�!!�V�E��a�� �k[Ҋ�
�!! "y#_W���vP��XKg�~��c�S����i�?��L��@�6�~7�C_#�D�J,�����p�I����11���(��77��^;G��ej9�.oac�q�Oh�QjwY��>,�6e?��U�a�x�?������\��4��LY����9ِ3u�W\��
#��1��%fo@��z��^���('��([���W$ץ����>��r�k�ܟ���9S������<.���<Z�ye���@�'�=�1�����p
�E�=�eLr �{%=ʵ����QXA�qփn��a�(B�D��nCFhx���
��T�w�J^f�I�3E��ة�wו)Ć�J������j<N���6�c����/�C�#>Iごm�9}O �|U��AC��Wk��j�0�:Qyt���Y���æ�3BΞwT���X�f����K���[�خ�����$^�^�a���]��Q��;��(�<Y��\�����:l�K��.�T��T�+���ּ��*�&X��'��{q����(�viu�AH�jY��[�k�3n��p�z�~�S�}��nԑ��QTB9n�b�"�O\xvA+�5Df��aC.?L��`Iü}pD��fR��L�@���L?�;T^f_�������:�΃�@�{sA�1F��B5}���o��Ӯ�J���qD�ۊ�#p5��K&�ցj��f�~�Hb��o1ʡheHz<--�����o�#{���?P�\۴|�	���tR�e�0���x�OD��B�@:L��H��/��^����%�}L�:�	�Wˁ''q>(Y�4,Zy�m
B)c���ҧ�X������Bew��ԃ�}���^�Zی�A�M�ȉ��P�����ݑ1�t=4�C���%}�;л����B8��~�����M��:��Ms̤��W;����'�n�Y���]a//��P�C]���Ɉ�S��V2����=5�sR��;�\��s�wT��ʗL��s���{��dE�.ތ�p��֊dF����hĈ�|.U��ډ=����,9�8�x��
