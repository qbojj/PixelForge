��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0
ܜa���@Q]81���,"�ff�a�`�����)�&��ɀ���wz���:��U��M�BC��9�iu" n�����7s��c^#yh?�{��<Fk�Q�V�ۖ��eu�6��P+^G܍�3����f�N J{%Ap8�<˚,��4F��D�Ƚ��+�@ar5��mPY�4g|�r2��45d���Պ��W��hxl'���S�-2u&��/����7��]�q��ZqO6���������������.��C	�������T�ȶ�p�W�je�]u�SG�͌���o:%��<%Y B`��U����z$1!pYM��W7��A��Λ.�.fy�w:����`ހ,N(@Au��zl����g�7P��ʹV3{�%gSt^ټ�j����C�xŸ�4Y�1���w�(!ƽ;�,]�k1��C�7#��	��z}8��9���,�F�|���5�le 9$�,fX���]X�OXA�� �t~)���R5xo�Y�I������%o"�$�h5���D`�Hz��3WܱV���/v�Jfl${�	��������%L3�)�tˊ�c��f��Hڬ�����h'�*��"�h@������"�e���%4\��.�U�2[u���5]��ĺ���5���FL B���{��td(�Z�~��H�;-n��z��ٵ�{߬� �I)��]▘Q�EA�t8��*L9�ٿk7@��Iuw;1�-��Ͽ<#�Z���$����ku��_���8\���}��\?��b��*�����JQh�v�����~��u�*�I,B`C�7|�PKp\�Y_BD�ȴk������K���H)����h$�7�� cW������c����Pb�39�SU`ٕ!W}�h'�)��|gb���R��KI��oD$����&��y�ԟ�2_��ycl"�j���^�z�Y��������|��m��Y+ߡ��j���ķ@'9p�Zܫ	2�,}��C�y����E�۞�2�0`Z�B���:�~��H��9���'M�i���@(qcE��l��
������Mhc��"�I*���j�.���4��蝘����*�J�ie�S������$Ѩ���_$�t>�4W*\���l��Y#ZZ�ޝ�}�}^*�y�k���̤/&�Ι�z��B;N��"�<�gw=z^�SJ���G=
�����tV�y����ho⁫/n�"�6���zhZʹ#���q��k�wXg�HWQ�{�X�䢴��ΡRJ��A�2�^�@���ɿ����a�oW�:&��Jk`O��>�S#iE�Ƃ���Ҫ�iT�Xv�n��9�mQ#5��oCs�J��{�{�p�P�w��7-O	�(p=�HvR��ɾ�ڞ��w#�t��^�z*L� D����pn+\�,�@M��[��XT^�ӭ��q�u�e�
�D;̡��J o��T�y.\k|�}��u$�L��V((ؑ��o=�� p�4�3Vڋn�l�|�ińn۾;�j8F5�_ԑ
��v��ȜO^���M:�����V*7��2N|���o�)������S̝i0��ܵ[#�'?���
����T�N�����J���C(ݾ���Z�q5Bz�M�0�ϋ�

y��K�Ϛ��ƐmS$�V��?!������ɍL�5�o���|���QW^���ɦ�+���{u{wZ�/Dnqu���GZݪ�0��Z���Z��OD����R��)1���wjO0i��k��|�/�!v����0w���'�"�
h$�s=�� ��9��}�2Ϳ�����e$io2=����G�������D��΄���c��Y_>��G��S�dɜ ���h�i�v��ݴ�&Dཐ,A���1.{�X������B:i��G+��n��Ţ�p�����
��U+� ��W���c!!��fG`oY������}�<����|l�5a���ޥ����3U�-����X1M���9�p��(]��A"�.����7��)��q�]Jbj,�\_V������#^N�l�x�G'> C�M��61^�I8C��L�ͭ�r���ʆ���i���c�bcI�{zx��#Oߐ�s��n���baOV~��#�O�$]��5�|�g�g���`�n%�G��ƻ�=�ᢄ����Q������'�Z�35����<C�r�tV���~��!6��4{F�=��w�}
Z��m�����#q]�鼷s&�ΰ��U�_.8��9�=�L�|���A�Aۓ��q��������J���F%Ok#��l�P��X<���O2⨊���������1������>��I�L��w�i��ְ��]"�\����-�G�o��7��MX�}F!�p�K��'�]���ڽ�\.]T7h�OҶ�B��x�� LlIUJ��2�uk��(�q//T����*���fD��Ox�6U�h����i9ҹw��?���.Ѱ�!�
 "�4��z��7(+�V6�q'o�oR�V�?�>�$�0��c�D�k�D�7�7�����y	{T�T vd�3ans�8���Ƞ%�\j�	X�X����@U��n���q�X3��W0���,4]��Me�9���~ٜ�4?l�yIw�կ:֝�+��e7�"�%�>�/Ry��R�S�@6������K�(������=�f�9-_�|�fl{���Ӝ�#������t_F%�&�����S���ɶ	4��`T1���Ə~l�E�G���CGF�A����c�=�P�p����V9�W������ہ�~���|P���%�u+�K!�����0� ��]��Q<����e��B���W��!�T���������6 ��"a?9	���N�A;��ㅮ	"�A��-P���R��������h/�k(�;L�|�����F��˜�޾�ښ�����k�����LE��0~�ٔ�	��]uc�?X�{��A��}�F�tC���Q�$���
����*�@���O-��5/���Kv#��b��fdb���9��ʮ�(��H�u��ԑ!u6����C�R��&��=�����ct��ʎ\�ga�E���`n�	X|a������Y�Xh���
����U�ez�!�*��5�����՜�bvH���JZݎ��GW	μ�Q���ֲV4�U���M"�L�V���+4k�v����g�"�Bb�����K̍�;v����k��TZ�kG�����0��]\n�x�]�i�s�E¦�U�����t���;+Vy�(�x�h�t�t+^�p@��zf�\x¥�
q��û�=�A�@i��$�BJ��O��g
��J[�=NۯB��e�[�Se�@H�fb>����[b���6h߀oV��,�*��8��it�ʏ; �5�}��U�JJ�҄�'ʿ�{�u>3\�ׁ���a ���PZq����g�sَ�6:��.�2�V9���͘�����39z����n��H��O�����>-�:T��j��Y/��o��Ӽ���	IjL^f��ޡw�E��G"_<���Mn�_	������۔_!� G�W�5��7�p���5L�ő٨���>��*!�:�����1���Ɇ�t5:m��f��� 웇���"���0������m��N�m��ϰ�����؀g�@F(�*�[v���i�	3�%�8k�p�K�����m���"��Vp����i���3q	��"������f���m��N�fg4E��G�_
W�OY0?K?�7���s��;�-�w~bNUGd�l�bў0;r�ȇWn��o�51JԽ� ���ּ\�Ȼ�p�&�_�x��M�j���g��2��F���K.��v�s`L�4��Gq��|3v���#>��B]mۼ2A���}a��2�d�6�5-��c���?!�q��ث_Zu�9J�f!��Z*�.`q{� �^��6�/����Z�.�/W�x�<ݸd�?���ٰ��
�f���1��V�6E�;����]&�^��S��(d���މ0�la��]Y���Ý�3�H�Q���mY>B'܁�H%G�.���)(��j�|fJ�$\IF/X�!05��{����5:��)U���1���"�sP�WFY���{�Y-�0_��z_�{{�*�V���u�<������[v�"�J�����u�ZRl�P!wNm��.�l�8A��--K���K�'��#W'�#,kML�5~ 1	�}��2����W)�נ<,�b�0��گ`�'��m݀v��P�2���1P���4e�������l��#���M����LW��1y��w<��| �`�Ӏ��R�4<���[� �R/����T���Auf��o����ۏ�slk'�5��D~����I?�Č�I���(k�dS�_Kc����X�ݷ���X�r~��X�L�cN������+�V��4�H&��A�Y����*y,�e����9�;��{h�?MX�~h#}�!.t3Yk����1�R6M&���
��O��z���=�%da�I-�X�{k�jo��f!D��
����J����PL?�4G,���7w�5�Ka��}4D_[).\�.v7���}]�?���M�0�rK+C��
I�nN5P3�����KèA�7�t�Ue���X���
�c$t1E������v������`�rW?b� ��艫/�r�������*z�{i�ۧZjǮ?���F��:�t���0�ŕnl�&��^��?D�x0j#��������/����z�PH�_��p&m��Վ�`'�`1�7ƾC��~�y�����v݅��,a����'�Hl�G��Ϝ)�.4�G6�L��yM8����χ܌�Z��;�jz8{k����<�ő4ڌ�ږ�T��m�,[�lkT�lj��N�g,lJaʂ,��
��$�{�A��`w�~�|"��e�鳻�ߢv77~0��>��TF�w�?Tks�?	�]�v�-WJ��g��X��=�D3���q7L�8�?�1�b?��W|��*sُ<���*�f�'�=E]nfN#�O���\�cH�*�kϝ�������Zp+�3-?Px\1�
sl��`�M�]S�Y�ޮ'�}EL����n��o_���tAt� �b���Y�7I��s�����ќ�`,��Q�5c��l%t�U���f�g�ԛ�ag���\3�y�d�k�(�����]��f1ڽ-4��/ �E��CI^CCi�(�T0�^�ۘ�o�����t������?q9�c�!�do�X��.�m�i�.�Lai���6��B��	�1���j��ܣ����%���]��I�~��aP%��=i�����/���z *n��N|�.3]d>T�/�>`A���X�>��d ���B��#��S醸�q��,a����;�37���k�Y_�T^�/��9$��Q(�zh�"s�Ď#T1�!_���ca�b��vm
����O����'��D�U�?�AG�%l��(c^��*�8�e�%@�v��>�=��f	np����1}�e�+�Vr��';K$�z��
U��7J� {�s\�|��l=c���l�����K����\��C��MXT����~���1�������.�S���J
b��U>����4����u�^��+�� "޵G =��.A�[�c1��@�xM3��,�1�n��9$	����37�}N,���Z�'����4�q\{lK%+����&A Y�����ꎻ@4:�\4�����%2C����)'V�,a�G7���BFU�6��1��n�!��v�G*Q3��-@�����Wi�V�ԅ���k���!b��J-��!e���S�'��:{��6
����iiG��bn��
�>�؂�0c��a�&��e�zׇ�_��aQlw��{�������½`4��y��Z��2�W����a��5V�^�1>��G�>��m������&�0����{����'K(�h�H��=�9�X�(�h�4��P�4�@{X<�Q��M��|��cWI��,��	��2�+�G�+����r�m�;VT	*�����k�K�>����&���^��9D�
&�Ӣ�=�HW���+5:H��[����+x��|���TH:<�J��[����ʪ�Jn"�U\��#>_�z[)s.��[�N���!u�g	�h*�x�qN�J��3�;U��sY����A��05ɇ��þ��	w�ڱ����ޅ%��/�7KQ�R��/�f�Q`����zg�G����`�j_�vp/@i�16T>ބ+W�dAr��n�K|��s�" 4�uq�j��}��7�K�� {�K{B�E�Bu���M*���P3�jD�#Ez��ޜ���Ͱ�]���ȉQ�SwBw�1Ot��C�`s�Xq���cAU�%u<���d��L�h���~�I$݌�Pu��}
�J��̜���yz��>��M����נ����b	��znT0���H�*M�����?M�#��eA���|�|�\|�O8P1y<%�E��pD:��@$�m�m�oS���B�,�W+�_+��4�'���Q,�;^��ut�q�7�PJ���2�Z�iƛ@�; A[v<n�[�vŶel�=,.�)��
��=:]��	�E�_#N����t�ɬ+��ކ� `�!@h�56ETz҃��J-Y4*Nd �u�g�� ��o�U��R�&}�$�/ܫSb�Ů[�߸���@���r	]G�!��!7]��c/����A�<D��GR�l�>��U`����n�[Ǉދ�P2O4�����CN�̅^=��br��q�� q^EW���&&����B��_ ;I����FFz�+����M�&p����^��n�1���7K��Yw��;Q�SZ�w�#vz�C�53 �дc/(�!_������9.�͆,�β!K��X?|������>O���'ح�;S�{:cx.F�)QA����CS�$$Mz�
��ӄ2W��D�٘��$N�*T�T6����nq(��Ғ�zE�����r� <���C��s���W(\�pBF�<�D9�>e�r���h��4m��%�4Hyu�e|6��f���_Y<��r/��f��Y��7~Y�{��t9��aa ��4l�8�es:�9A�?��r���'�Z������!ݑ��v���UCF2�厇1��͛Y�,-%H�� �� 3����ai���򙲧��m�����N��V� 9�l�œ^>Ap`��u撜j0�m�6r��b@��/SwZ��k�[E\Ѱ�qt�>�Cᶌ�w���Cs7:[���?;άt�7�Ih����0�����3��qӣ���\#gm@F^+"m
��=��AMt:	�g�0mK�u������̳�MhkS�(Bnٚ��?O���I����[��q̃�A��aھs�p��������P��">E�R�a��s���A��h����c��sq����$^��˾5%7����}�!�AB�����9�,���k7�K�ɰ��9K.�BEgjH��m	����pmCDg7\r�����f/׍�T7U�����<2<{�!�~�K>w��~���կ�#nd�B��S�8��^�H��;�g~�o�G���� �^ѩ�JR�u��>��8���bA�}���V`�v)s�������ّ|��Z/��s��4���i���ͭ%����z�J4W�;�8���8ڡsȈ�&���0�PkKё����`��x5����O�v�N�٬�)�-,�j`�}�2�H*�i�_��"�<��4�.6tlPIr�6�`�u��6�XJi�H��f��*�dMf��T����^���(�]�,�~&�x�,�5��/e�X�WOd�|y:�r�&)�* GCpz�v�����*���7`�	���29k :��b�+)����tتU�1���،�y����T�o⼦T�͈�o{x�����Gc�	?4�'���r��t<��܋�T�!��:/�En��m�����`�=C��Y�H��Z猧��ߞ�-%W!Y�WN�2/���^������q4V�a�\��U�F�H�&��X[7 mv�i>�a�
�~�lx�c����u)�zF2����|��j���p�ț�2e^�9�T��0V�?n�k������%���#��*���I�#�'�^�yͨ͠�9Gkb�9(�j���w+�e9�_EpJ�Sy������w�v�͟Պ��rUT����x�%�zO�?�����^]��^=O�P�%�;�$6�)n1��;���������_� o��$�5
�+T� ��7U�u�t9ר_�
IZ��K>��7�o�+�	������mkh�]�;��H�,�����oU��0��9�"�S..�/^��_��9�CIɢ��ZhW�/�7PΌ�E�в!�7�ʫ��������������k���E��z���g*+0����8�@]�6��v^�D�?9��r�������>8"�_�-9�i3�8̌�6�Zg%���.A�;� ɀҪ{���l�+]�Q�;� �����Rg��=U2�hi�����82�9a3=��˙���߯p�/���.X��P��_ފEU�p��D�BHw��aV�ѓ��E:��V���
�)�?�,�Z����0GfY����Byn�<^���	��7޺��y/|��4��?M����z��몸A�D�G�2�ck��o���xڑxb�3Csoݰ{G/�V%��\��z�	��Y��<>�@1#WOP�5'��]%���w����"Zճ�qq�C��XEU��g�� S����m�$>����6�����*��4V���%�C�їB`�â�[#���7̝l��~��,���ڔݦ�,Ҥ�Y����9�����@�=��9�D\��8�g(����r2F��^��MԞ���������
f���s_f��xN_vN��	mL���-�j�&B��AsQ�:#�~tEO���T�Y" PB+�!ܸ����I�[w�%�&N3��E��,�ʱ�Y���[�U��$~���d�~�Iza;%�׺��ai�����ǐ�ױ�5���m�z��}iJ�Qw�Ѝ� �@���e�j�cB3ta�yH�5D�qւ6�FL�Í-���:�/
ww�O�M%���0;���K0%�g��&�b���PR�3�ńF���&�՜彋,ŷ>];��]�b�!*�ܘ���<5�6�C�Bʁ��f'��N�h�/>�ēZ�UD7�560Ї�3�#$g��,U�Ʈ|XY/��l����{���3�9X�[h}���"��{�X��^�XG��,f�
y���� �ԅcL��F���qp�5��ڴ@�E#��#`��z~7p�B���Y9;��<�4�l4��m�Y�\�\;� T�nC�x<��z���ao��J/�e�_ ����岐9MP�Ԅ�s�Z�����c,�I�t��zK���LZM��7j7
���L����%5�;}��B��-0AU*����V7j���稘�\*�2b膹���ϭ����B����j��[vR�F�� �\�/�+��k��RZ����h�?Wmg\m�� �2�\7EƑ�]D�~=��Yh.��'�I�}�W��b��@�fCn`s�G��|lvӷ�yW��m��!4�Y>�']�'��Ȑ�uNқpMxU��۸���p6}�\4�X�YYx�-��]~Yգ��|Et#��e�K�$s�r�)� 7�r��A�)�S�ui4�)�|���گzחܩn�I$��	�*�#;�����e��ٌgR�?�T�����&���*����k����V���A��[]U�cr��ґ]�Ǣ�R8�����9���j�p�B���%�5�����qn���P��J[ �7���S��ûK]+n�h0v>;��XR��xݙ�JZo�2��N���C�����]��4���Ι-���H�#�E�I��r@�m<Ͽi�uٟ����S�:(�>ș�ɖ�&����8�j��U���M3�c7����)��AF��ҴQJou�v�3�r���Cfz�Q���!�֦��J�l47!J#�h}:�,x�Ox��&�{���E�{m�	L	�k�؈_LM� O��z~�Ҍ4���*�@5]�hW:�WbS�N4�9��R��������]�2��	6��#��/�q�"��[�����:���^��Ç㙒U�-hb�8���P ��n�,��$A�H�"��Z�)���:(��T��>��e��R�ل����!@�%?�/���Jܱ�F��'��r�݊Í��j��C{�+	<^��qUx�H�C�v�Fz?�"��$a)�+B����!g��b��q	#}F�G��b���2���iI�)�=�R�M1���������Dj�U(������դ)�۷W4?tf��:�����~ː�fO��\��٘�z_��4�O>MZ��]A~=��NV)a9���������W�r��b���5�:���g���[��7l�������e8��
�s9��WD#rZt�C^�e���8Ө�z95`7�!��d7cG�!��A���ꕙH��uc�%e��əw��򉢺<9�fx8Ivա�N�A�����!������]K� "�6;�%Ќ`/E5��E����G�����&������,Fh��.Làc{�u�j��0�Z������g�{p9/a�pw����gV�,�ɩ;G�sk��@oj��PG]Ǐp#�g+v���nd��?����R~J�p1�:?�)�w��0gd�S��m|\s/� LB~��Ϲ���\b�\�yZ*0|ڨ�[��X�(�x2�X�V|��f��V�(�4��F����S�Y7Ĵ�s	�b�ҝJC��O`�� o.X�f����W���	�"8�7Y�jo}�NByu)��z(���f�-n�̼���˾��eʈ��\�"԰�=��1�<�������_%ߥ)j�p�}l���@<�%~߷��2N�����4[�(c��F�s9[�Ӟ&��o.>zUl���,jl�1�oCY]�fG��5|��B�KЉ��娫��%�bN�w>
npev�9��`3��֦4-���'ːs��E�t�*�}x�T��7�w4~*8��s-�ғ2iHd����r�E\Gpą}D�m�^��op�ݔ3��%�v߅'|�v􏍮@���'��HTq�6]����<����]T�Z{�U5�pH����(#�5�B�ͧɇ�L+���M^
~/��Z�h��N�`a+���J��y�Y(�Ot�N��lbb�i�j8���1�^�<�0
�����R�H��<��-C)���'�����V�Ȓ�j#��0]mm�'�^�x�Y�P��y7�aIR�M��V#ϨPDh��ŀl�����E��P��ۣ������y��"
�'f��O�0W4�4t�@\�p��c�}�
�-�h��N����m�\�j�V0x�r_�ldyV���n�q�(Y҃�\8%�-r�q݅�H6���+����6�c�p��Q`��?d����p^�n��Gr�x�tI�aF���n�7�B~.I�\MbS�pf{���TM8j,٨�Ko���J�nQ�ۜ��ܷ�|�^������b��t�Q�_�@��_����}KoMv� ��v����f��P#�TQ�.�!2Y�Qj3��G!��	����i��h|E$
�97#[ 1�i���d�4������ɴ�#�i��p�̻�-�?�۹�,~��k1���q̓D~�l�����Jܷ�ԠEX�Ȩ7�E3TDL��X��P}U��k$0H��M�C�GX����W��X4����e8�г��C(r�bTQ�f%e��2�t�K͌#� ����rW�A��*ӹ7�ܸ9��<��\��u���>BEމh8�ƨ�Ew�>hW}� ��޸����Na�����aY-֘��*��Q:�o�i��y��d�6�b1��7:���6�;�H��Mۍ�=��?������׉���L������ IR9���p����6�j��������N�����-�E�Ny����(���w��>tF����1��:�g�PI�Wҫ�M'v>�(��}�Ν��9y�X�V�q��Y�f7���e_�lFѩxJ@ 47�m|4�Fa�k(�0���"��s���Ю�Vn�^a�Ǳ���C�I�}ߛ����p>|��
���``+/2h���.M�%��׆������5���<q����dZA�@�AN�Y��گ�݁Y�����0�Qc(܊��>#e@>�-�(/�U�u�P�����*Eܹ^NǏ߬�%�o����nM�f	�n�tכ�u#��ׯ�(Ҹ�:M���u �,�1*V27�Az�g�!��XG����ՙ�w��+���Xg�)��۶���5�8�щ�]��ip�cw�:�Y?)S.Y�(�L�����fe̠���e�G`�A:��|�4¬2���=5�N�h_����=ӹ�2�T�R&z����Ѕ�_� k�4�{�R��jw���@���M������Is��M��c<s�pb��-���
�ыH�QI��צJٷ)���^Qi�ﬧ:��i9�l�u`m8��IY���T?�A[�C�VH�U�nv �'��^L�,�2���∕�	QMJG��&{d�4�m���a�\�Ƕ�&D�%B��Lf���i�ĈEG�N;��K3�V٬�&i���RTR�����+� T�ڢ��q�:���B��hE>���XOl�a���(��f޸2���c$H�e��_����*�C/ҍ_�f�@|b�`v��WL��5�^���r�`�8{�]E���ZR����JȅO0&d�`��3zAs������ema�)' .��x.�>]�_����kq��~����@�{$��c6�?��t�h��Tg�zV�xC!�����k'�..����|Z���SgL�Kt�5h(5�Cr��8��A���\AF;"���]`��7�ճM�1��T��r�P�1=������ڑ�v��k�)��2�Ǹ��sUW�k�#I%OgDxܕp ��2�п������F��ʡ��>�����D�r��,F6�=a.L�Y��ju�^����y};�K�'�fy�&�_�<Jx����v����FB&��*sq�U�dDXYs|{@�����Y�������F�W67�w�*�U��h�	��AfL3�ٴ�ю֯W>�Jgd0`���<�3��)�X6#�$�sث������X��&N�,5/� ��p��?
~U�W��e��S�����3�q ����-��b9��b1��똄s@l�;ٌ���H������ď��ļ��tEI�c%C��T7�y��s{N�5�VC^+Zn��\M��E:Z�l`�V�^��[�!�UQ`�@�a��m�J�?�sN�0ﲹ��9�O�������D����"���J�d�'��U�A��#�j��騶�)���2���ڧ�eq�,��iޱi��<����G�������F7'=�	1�/�,)B�.|8y|+��ʈ�Mf0;g��H���o7. G��l&SxEK{;��R�`{S�
z�h���a,�V�҅��k/�E�ϫM
