��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���pE�KWvSj�(�1,�^n����6�^�!�A-(ΟZQ�����S��J(ִ)��t(�E���:v��u���3���գ���URO{3;}��l aI�B�F�Rr鈇hI����{=,����K*A���y��kcg{�;�d����ف�m���F%�����#�QN�+���G0�f�����x�0y�Ѣ��<��D&�7Nj�Yx����(���{�x�3�h��&�#��h`��6�\zm�y���5�/�Y�:��roAG[�L�Ϲ��e�Ӭ�џ��S�`Y@r��� �K/�\�ʅ8Vf��_Qڌq{Z�k�	�,�����E����KD���a9k<��G>v��U=
Ɋ4��k��&[#@��F��P�K�xC
�����̄��&���7 0�a�zc���R�ϓ ���Xw<2P �l�ޙ���c+�Wt����M<��W?�69d�	fʳNv݂*2 .�5˘�H�L�9��(���$5R�}�y�̜{��N{s��a6�l_�Y�}�3{����S�� dBK=�n�B�`��ou`������T�Of=�3�T+��֐�ukӵES���a:��IN���Mw�A⌺�wK�D�|�F���b�j
�|q��5P�[������|�P��A��W�&��V�x�.=d�(�0�?�=ȕl��?��g���O3��O�1Y���4?��p�1SEt��}R,S+����?��)�"T�t3O���ЀӶ�ʚ@�H~��s3���1b�h���Jp��Q��o��d^��	0�9,���mb
el���T��er���R�)�hyM��/0���h4��J���%fGM��+'���84ͬ�f�JE�z�'�d��r^��+jp�8_���3��S�W����.pu�X���<Kc���J��k9Թ�(�5�����VK�� �n����l{��I�$ʜ��ma/���G��hY�P.G�/�e��]�'A_��m�ͩ�t0�9�P�W�,4���^l�gmFQ_t6�A���������T�--���gS'�L�!q�M�1�ţ�������
�[��0�ܣlхE!�o`s���������p8k�PQ�&qr���c��<��n���41�1i1���,Qy�oE$��������UE;$DG)���׾o��I0��k6w�YH�"X���__b\rvu]���S4Fd1���fYS�P��f�ȯ�:?�ѬfH�������͘�Z�1⨩�{87+eZ>)#��d��yӔf�y���9/'�\��!�S�j\����0�\b�a��I]=!pob@
����e�I�	+K> OS��-�r������}�w8Q�r��u3�W�6%�}e��DG �ClO���쎨P����/�vᯯ�*�1����n�~�Gm<�e��Ӣ���d4D���jE��d��괔����$�+S�{�I�O�hz�E��x�r��k�p^�B�6[����]k��;��-r��ˀh��;HX^�X��n15_oM\C�B��0m?4D�����}���Y��^؃��,�"�vT��k����FKmz�㛵�-C'yi�13&�樬��*�80l����Ön؀S�g����I!R�q��5��r�
'4�h�g�X�e���*�.�fH�!Rׯ�_�V ������d�����4�9��< ��P`�8og�C�7$���<W���2ZHrل\���F��~�計��)[/�����V)�+G�*���5�1o :�]��NuC�4K����k�&�T����{	T��9w��uZ�P����h��4��#0?jQt[�� ڏ��pMniH�=��4�ʽ���Qpq�(꿙�ɋo���ɍ��[�̜�VOi��XAP`r �<���#�w���,�܆o,FE�<,y,��Jm����zo<�P��cϥf�H���߬��Y��
�B�X�r��>���B�Z�<�U=�֝� �0��3P0<Oa�s)tK�ACT!r��mv`)���R̴!�9�|��`�VgG5���1OK�قW���T��ۡ3�	1��)>���̴�P��8}ے���k�$Y/Ӆ�d[{K�+4�pt��U�߯@f�����kz�╻��6d�ˇ�7�=c.1�A�L�@K��j����Pk*|�5xV�7� ]!��(6OǷ(&�ɑ%z��D�т���g�y@>���*��_��\5c�D���D�D|H	��u������EV㝟
"�doؽsf������|� L��O3!h��f0ʗ�����R��KD8�
L�d�Pч�By��� 2z��j,� �77���A��@b�zY�4���~��P^�t���'ҕÖ��H�uh�o~YÎ��ks��q,��x������Ώf��	΄��*a��2CN;+�^��d#�(e�J���׆�j��Մ%(1f�D�hĒ�t5׭VeI���4y��Ħ9c���7<X�t��(ExnP��>�漌��U(�h�]�cw_��� h�O���pΝQ���evX��'���OS��ߍ �'ěx����W����c��=Ƶ���iO���3F�=E�9��t�11�xxG3+�l2���;�r��H�0ٙ��[��x���6P�$��&���5.~��l�,�� ;V�0��-�u:5z���<襄�r�A?RK^�L�4y�pvQ�v��\/�'��E)矅/c��Tl�N��a���.d� ])�h�^����di
�6�έ�@�:橏��t����]dWX���<�u�m<��%�x]�5D�b�}��{�W���K���pǃ�,G��O��g�C����-~�D���!"_s�H_�^,�Z�19$F����3�w�tK�M��FX�X�� 8Vt����.l)�����`��>͓(�ub+�~�_��<�x��#�r'_'O$�u�[�(H=�����8��)^���(�U;�ݜ�Fg����3F��x]f�Ѿ���t�xn�q���*Yu?v� �a��-����J�d���-Pҝ�-x��ɲL���	�Ze9��I�'�ѩ ��Tz;LuA����8�yIn�];�4>�;k�t���p/�rg���ZB���-c��)������R5��0���Qm�SI�n��ݩ�Z�'�{���N��X��	�3E��}a*�����CW��9��W?��m����u^	j)[O����&1�H߀���R,�J���U@�N/���p��~����t~���:��j��� Fs>�@���� WO��0,����yW�ސ����� �(+�>xԮf��)$;u\����E᝟�v�|P��g��U��> N�B�L�Ҝ���&�T�x�@��}��zXfC@-���b����!h��u��;���x�O���笈c��J��F��#(M�<5�m琍hu�]�
��/�82��d���l�!x]����*�`Z�m'(G�ڙ0���,�@�x��7@	��>�zyY\��T�	�R��p��j[�J*_ګ���b
t���l�~�5!R�1^X�z7��3c���ȼn�6!�I��T�j�Ɖ ߾%��L&��y-[��&�+Y���;,�o5���0���t�2Ri���������� ��� �@�9 )�t��N��m����]]j�{b1(�LI��*Y��*N�}| ��<��V�x��3�ɚM��p��<�	�e(��f���܍�0

^�x����Z_��¬��ι��IԈ��|��X 5�c�"hKD��u�����2i�F���D�J�6h����f4�{0@g����(�<̮>����% �I|�*y}���ʌ-y�h]Q��+���B�,�Gjû�q�J��tY�)���f����H�EQ�8fQHw��IK�Q�����&�v�/�������@�?�ԓ���`�?�k�{1ׄ\s�bu�^Q��P�գ�V?{�	}X��ʎ��A��iF\� v���[��'؄o|�q��b_�pL}ҟ�1�n�+��虨����|�P-����e�q�Vj�������18�ǵ�T�!���}o?�N�KcW�j��v��(�*����J���-�	����gŊB~�+c�rZ�R���ń	$d��0a1��X_:W��҇ԣ�9��гG%8�����+/xc��i�<QQ�-�\��VGBZTrP��u�.Nh��cVنl2�)?���dG���ݮ|�c��g�m9�J�sU=���(����Bs��)2�`����l�/;��c!6��4޳�Q��-hќ�����N89	���b ����OW@�d�c�|��Ca��S���m-�ް#<ǟw�쯫QM�^ϜE�Q�`���3;u훀9ј��]r��\�AJu�P-6��(��b�,L�/z�sW[�"�<,U܁�Q3�Y�C���0����7BH�b��4��P�7�%i���~�Y�1꘻�K$���o��ֈj� {�S���0���0�Uz���1wy�$��H���HO��g���Cձ�.�1�̾��Ni�%��S6fN��CQ�C$�����9���a't	�e�$�1���,�j�?1�N􉍘�=���Q4ۋ��K��F4��fn�>�m��6�1eC�o��1f��hƷT[��s��������5�����e��:2����)��P���Z���&bL������j�&�9]��vp��)Ti���+��59��v�cm�&��s ^�`�|$�7���)؉|���@�5���ߐ��՚����ixW��[��K�tMhw;Kd:6iS��d��5a�7諒&���4��*?�Y��AS[���a���P��5�f\ެP���u^ۢ�&c����/�-
)��)b��TЊ�j�9=#7<�@_Д'��$��*lC:�/pE���ߢY*3�� ^����~G�cx	q��	n�����F���$o�ܽ6��}���n�% w�F	�R�_��.����[࠲"�ޫ���O-�c�AF;OA"[eWK#�l/�+,|���aRx��D໪H;XR�N/̻c�a�~}彙1����Q�''b�.�ѺX!#@<�,�Y���23a��	_e�MJw
NI���8j��M�
�#�P�
М��ύ�)R
��7i�Se)`_�,��B5M�,;��ŨD�z�H�0>�ȁ��R��|ܮc�-3#r5m�"�|�[e����2�ou�%]��r��k��y�MW����ߡe�痪.��;KT�g2t��9�=�ǋ���v�-�|�X��7��1-�?n��"{��箒�rb�oI��%���r[j� '���~�=�.k�7��ɑ����N� M.!�1� �@}]�4+�0�i�MϻM�O�W�L����a��Qk��P�~�����	�����!�A�c�DcdZ��Jh��r���p};2�W��9�b��	�)�Y���+
h��&t�K�L������Q�0����J'D5�TJ{��q�zT�q�nA�[� 6�	��R�����9�~��r�"�$Dׇ���[��'ޏ���թ�ݓ��9�!��]ǏK�w�l}�[nPïw�� L���R���X/tc���D�&�.T�3����%�l���φ�/�[���~*[�˛��������6S !�f]��g�9���e�%�;*'Ó.�S@p;��z�4;�N��B�L�f����/!�u�w$���6�<\������Z���V�P�M+ &P�ʅ�*��k{^Gi�I�L2�H�l�#Bې���3�ʉR5��gq˸$��n)�ܝ��2ӌ(Gn��2އ+>��8���AKʴ�?X�Dg ~I��g���`r��d��u��4%���"��D82"�_p�b�&��W5�+�MG�鉙�npZ+�{ӆ�`�Wr���q�� �T�œN�tM(����v5DO ��+*��^zH�f��Jfu��1�
