��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�06���A���ZK��UW��BݛG�=`Ŗɷ����ݯ�m>�	,P��	� ݨ[~Y7��|v���lp8{^vc���c#7���L�N}� �"WZ-�vɲcL�#�|���G}�\r)�c#�@=�;�lM/jr}r�}n�U�LxF����[?	Ӛ8��9H�� 睭�8�{Lokb�jz��f�7}c�/'�@A!���{�:m�� �?�H� ��fza����§2"���S��G"�v���m��h,A>�#NnN�i1���!��:B��O���K30jYǠ�?�EN]iް��R�o��nYP_�#a�]��-Ci�a��i���87�~e�@���c d����f�80�$��H�ܤ��є��EBV4x�&�5O�0Q>�3%�W70�с~F����Do�YT�Z��z��̈́Y���ܓ�|O�����#2�'��!�ڻ"pb�P���ZC:����y2g3,�^��W�vz�����yhIf��w&�2��<�M��l�G��7�GmR�cScj��ZBb���x�b5�~ ^�}'<-Y�9l8-�S{�L$����_�[���V�2{ˍp�j��r��R�+��Is���a8����ct
�;4���[�ԁ*ߢK5QZj�/�����o�dKA�L����3�:5z��GT^����b[�L^�����󽟙�He)�d�#�E�"��� ����/AG����D-B��K�!��z`[>�)S�%ߪ��K%��_D)^��I��ҶN"�*�@���;�,�km�F?�|=Jv���H�p����;rS��N1�*�Ac�<�����]4&�lН5bF8��İB��~0"N�Q�����3�VdKb�
f�]օ�ڇ_�	��aWs$�]1J�6�`v��}����~JJ�f���l��"�F��O߲�G3Ʃr��qH%c�ː�i�ꝋB��	������m�f�P�)�'��k�5mB�{��=QW�5�(_!�!-��U�g]�ng��'�b��m䀣Wj�D�%���_,��������	)��rA��jt��J��Ί
��\k?�9�V�3�9���Ee
�ʲAn�7#�=�\h�>JX)�H'")��80�)~Q ZM�*!DP��˴d���O~�"��^�/��I���>w;�lY�������N^����x�g��um��M�֪5bG���#�{*b�c�ro� (T�(ƣ�&�ư0sp�_/� ��B��\u�Z����wPx��a!m��,O⧜��/eGq|9��4gʠ������ �l��r�+un[���s�~|�S��aN]+z�8D٩���g���"K�0����,���x���(�2^)ì��I��>�KC��-u����q w�%+L	�9�L�rnDSi�˥"�T	�g9���&���6k���'��o̴bl���T.���l�0�zg�}�2/�m�C_�o�Q�+�-�ΙDj�F;i��+�j%1�q���w^2�\g&	v�^��tK�s����>L0��υB��K׊' Q�:�v��Z�F0�/Q���5�z����c�?:��}j�ϛ�ٳ��ϊ%ɖ^o���d	��m%�>�U�Έ�V'����������<g����|pW���R�Y�=-�r�ê��"*��j?��>`S5�;��%�Y	Lk��q�-�$�`0�xcz&� ;���֦�l�Y5��>tzp!�G�gk�UHj,�t��C�J��6�t$ܪ'�'�)��ՂC�� @#�m�OM��� �R?b��Fq��Bv�A��zF�4u[_}�cwf�~�Ky�h+��tF],g�À& d�:��}#f=S~x^=�W����`����JU\�#,�>��̇9����^����J�c���Ϝ���7�<����E4�v ��
�=��zfAך[:��b�~�q�����Cmhaz�h��D�\��I������2��̻�9�Gl��9�����"9f�m(J��&� ��L�W2C�4��s/��Qm���?5�Z�����PC�;���V�v@;��mw��]g+�HY��A_��?*�� @�gq"Y��7R&7�Sx��ݬ����PD�k���� ^��
`;vc_���IN�kp���<����r�]K
�+�-(
