��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��sa^s����Hw�9��≣�Z�T��9��p34]�����4�N�9��
A�+j@"a���sI�^��<��5�04���ALc�bl����t᜘���NRјURf�hy��\�q0����C��_HJP�Ը����/܏�xT�A�> ;�!��l��ȃp�)j=�e��7L?�<�����s���|.L­�����p>eҫ!��B���z��b�Id9��5u���E�>��	���K�H^�� {�& FR����_�����h��睇a0�Zd_y�`��q�$��q�C���jI�5iz�g������m��]�di2yc<��@Q���@:��e�y%zk����Ё&��KY'l�-�[-�)G$ �KK��T�H�]�&���\cܼ\;87��d��!���	/���W�HC��_}/�Ͻ�h�����><�r;���l��-�}Gw̆4M��']�(�ޥV��~�3�5�)5HM� p�GL�Ȅ)��n����e^��
���TĿ؍���
�b�~�=�C�*QNxѢE"I6���X8����%���F�D:�S������6�F4d�A����R��U�>���ѽ�Ԍ���_}�ӓ���U=�X�t1���̄t���x���Q������"�.J���������
�-����u�=���aY��u����P�Y��M��,���;��(NAN��6�`�
�Tqܕ�K����2��b���.m�W�+�#�W�(^|�]��9�R�R���:S��~�2�d��kUʑT>�O[b� x����.�<n ��7�ȡJa#>�~E�SO�ƶ�V��"о;m��Ė�����a9
�D`�Em�^����2���%پ��[M@���T,�W�44vg�`��o�g�j4�um~�a�R(����2�gԀ�j;an���(�@p�\B�����qF���F�>���&a5U��h���&:�@�/�[����z�o���d�����Gfe6�z?d�a4�:�@��"�v�XnxG������+�2�A)�I�aҖK�{"��.��l6����YZ�6}t��)�x�.�f�v-���ܪ� �N���%(��z컢���=]͢��1��>[��y�[�&�.���v�F45*�fk0�m����4���PvPF�l~�	6aoQ�0��	q:S��XG2H���[f�"}�5�I71��"h.g{P�w0��5����F8���6աi��.R��N����)���c�24G�$�]���S�	r�M�YA�B���4�O[���*���}ƹ��g��Jg-㗭��;��9l}�W��<�:��뢎KA��S#>�9B7mRL˗2�����@,�D�G�ged�Ns{$�Z�k��u�L�i�����y�6����S��0'�i� �W)X��i�:
�iW�-[ͧ7��2��0����,��i �웥D���9\z�"s�.4+�]��1n3R�`�e�i>����`Cy}���LJ�/�f�K�"����T����.A)���c"����W��[Jm��|�N�$�p�����; ��dX� <oR���,é2rڞs/�9���ՄL�Y�!5�5�k�
X�_��������iO�@rD�X�Q��T8Lgt�P������H_�T��+��(���Ok2�����jݯ��E��PI� �&}�xs׷�r�tf�5z�L�ݏi����.�E�Y+�8���Xo�^�a�tGA$���c ��ee�GT��b�e{���+M�t��2�_q�@"��e5����'
���S��L!�s��N+����N�Ps��*r�mN?#����i�Y�	���a�<�f?4�1��㡻Q�n�_/�
��`b�T�MVs+lP�^ɍ@� �i���W� Ԡ
F���Da�uU�;k�[l��!��g״f�<�3c+7�ׅ)
Џ���e����;7;AR��N�7׶�Ӏqc⴪d����]���C9N�-o�a���ZP����-xȞ5����k��Ѕ�ӹ$uĵ�{�s�*�.�2`�---u/�F��
�Mp���_�-b�n90�k��W�="?�[��a^�]k�?*�o��6� I~Q9��7�'F�RQ����\�J��ň�D�@?�o�㔵�c�_����*+�DW�#�s�)����F*%���$���NnZJW�O�b�9z������o�����׮{�%C��Iϵ߂�j�>�O����ΉZ@8�as���#GUDp���Y�+ ��6kqϩ�>�� &dl#r��!��HPn��J?hGJח�EL���]W�c"*._��y��Ġ\y���6����z�7��|D��/�V��>�ࡍBmS�T�X��䵆p߄�YV[�c��`iܱc繐�e�{e�V!t ��Vp �}X(�'�;����W�:_��=�!���"���?��I��*�ݛ�Li���=KP��w�� ܈j��Gj����KF�KI���ءQ����Jp�4�o��(�S��Sl�"��]:!�C�I��qO�4W��������� p�I����oz�`�n���pK���-џ)V�
�ϙ�����S߼��������d(8���<�e��n�#.0���$��l���L`���W@���21CG���&т��2�����S����=�j�����΢݌��<t\�H��
h� 5p"�WÆ����K�����|jr~ي��2��۱d�tHTZ��N���$��6ֳH���Ӫ���y5a���TV��ݡf 4�~�pju�����W���<J�h,���2�-e	��RÌ����~8:Ch�����dǺ�1�*�k��ܖ3�y
�?.��e}z�^a.���<����f��Q�ZCi�@��5&5>��r����Y�d��,���1Ze�WKpi�am��Њ�q|����� �85샶����f@���L�r������f&
�ʣ���3+$Y�D�������ওhj�n�������t�@�1�v
ܛ��st�ӡD�i.÷/��֙OLs{�?����el�y!�&H������=���)bz[��7>�[.��}Ѧ�|�=����a���Ox��
���)ֶC�v|t��SZ ά�"��i�Prtjk��Ρ��
0B��} ,V��}�/������B��V�/aI�T�$���r����������q��%�çJ�\л	�Z1�f��>|,.������\!R��S���CMT~�ܠ�ѭ]����K�>�!!r�������yKߣ<�%7�̃��ڥ,?�T	��T��i�~֡\�Ki����M�X�����Z��=�.됣F���H�mL�B!>��?F�������3�vlK�ĉ�����E�p|Q���sz�ᮕ�ͭ��i��D,.�~�������8cw��b���[V���0�/E�ߜ�����#]d�R�-�����Q��	�Ο�b`���L�#� rf4/P�r��)�7?�k�&;���~��$�q��uZ 8���.�����JG��G�� p�,c��^��Z�G3	s#f�%�Ԑ��ࡈ�s�w]�Z01
�?^�e��}��`��PL/͡,,�Q�o~�Z��7��]h�%ʅ]��Gy=#W*K�JO��w`����jDe��2P�:�'L�5"�hm�j���Z�ǳ�����7�_��ξ���-�P�TU@�����i�-�)"�|����xȴ�
n%O7
kc�@+�#�����!|t�M����:h��8���g����+gHy;���~��ՉgDi���f-EZG���݅֝TN^si��q�;@����,A�6r�bS�0c�OEY��ņM_SF��A�ܱM(��P�	���������)^^�!�)��Ea����sQ3d��(���#�)� +�f��y�0.�B�g�(��,	"&!�n�L	�67??�\[.%r�ҧ�s6�H�����_2��i� .Ѱ`\����Y���U��8T�m2+����'g�d!�J�B��F���:�R_2�4<ܕ6%�x���7k�ut��c�f�:�6d��ڞ�"�4�����΃��Bٟ�	�_K=����ċ�:��J��ΉK�)�-�m}_�᥏������_5K��F��*��N��O�"[�{أ�kT�+��=�.��;u�}x��a�S�?��?���*qQ`��u�{�1��0�t6���n�)	�����65$WT㧩�v��7��x�ʯ6}��
�Q��I7���;�n����R�ٮh��5�0�^,ȇ�я8���t�w{�6_ ��CB��q��F�F�=ASgX`	-jI|Y��?��m�O
��H����f8F���6<��Q�yҨP?���8' (c=wN!f@Ǌu:�(��h$
�W���<\�,�Q�s�_o~A[w���5~xz'���h \����m��#%�ýU�H�#l����;�X��/�"�MZ�K��N�hH�Mlxn���VG�%���;O]���J�H�Y���h�0}�z
��Q@��vͅ�|����0����n��>�+��۳��P�������@�z�h�6��r͗������$p9�S��+i�]�-Igl�?��/�z�x=�@:�}lpC�M5��:p	��]�L�X�؊r���s���@��Y�G�Lcj��U���g��&]���B�E��pQK�#Z�������.���Z���D�E���"�z�rd5ݼ�ڀu=�s�Xry�&�Lc��	��O@C"��O�.�UcO;�g��8�*�0��\[�C{j�����~�,���z��]�R���uI��h���)�K��dm�%�OBx��.��O�*��2=�Gl�wS�~��6	bV��9�Hǂ�N�ƕx�žu�SW�Om�wP<�tB*��Z�X��́K��t ���f>�-�+Y�~��L�yH���.��0���{��
2V�i��������pL��
�0Ȟ�� ����J�������}�ٗ_���Dn���,I%�W���h�ix�b�ĊakQ݊��x��r#'u��ZHP�P�1G�$�qo���x��] �7��ª�Q�����nj]���<����ܞ�P�.�<A;�e����"�R>���v�r����ɡ�����~+}h	5r�z������8Ώ��\�5���Sp����� ^��L��~���UA�z��Y&�;[�� wz"iV���B$�-�=ig��`*98[f#�V����;T0v��: �17�jR�~�]��!tŠ���1i��O4,��������o�EI\���1�����Z�j̯d�YDG�B�3!ΝY�ħ�$��8����rA/;ƃ����@�}��W���F�/?�?H��{#��h��'m��I�s���l胒���r��#�R.��F����x�ү@� $�8���L+�f�CJ���
?Qr��s>ʵN̦�mO�L�i���vlR)��zhhXv���A?Q)[YP��3Y�r�Bل8�:��駡�Bӭk-v�j}@�!1�g��U�3H���̠��4۟kw��b)J?��Jl�W�nE�>b5m��N#�C��c�Kq����zD"�M�K�ße���D��Y;&=XA������#����98�}Tq�5|�~��ꊍ�����_nQ����B5dɲ])�>6tw2/���^�R���ق�z�G{^T�M�?*�YF5*z�wHխM���CH)���~�r�rt�_i�2�lK�������Ϛ&Pe�Y6�[�j$�ۃJJ����E�g���H�k�> ���\�FG��U�/��Mn)�3������b�g)74Fs����}�8�F�i*��WE<L¾.z����J�Z:F�Pq�i}(Ljtɐm3���9H�_�/Ԩ�h�b[�V�9�KɈ:�o��q����Y�n�ŧ�9�6���[!��?t�a�hE�<�	�2�_&nƶ�38�����}`�6?R����z���-騈���+�;�3M������Я%�,�e�Ņ7�m�]�SUN���T(��Pq�P�Ȭ͊:�*��l��h~fo������$2��,кJ=94 ��p���ۊj��':�/?(
K�t�E>8�-s/C�x'�
~*����C�l"[���~}�/'�xhʰ�?�C�Өg���A!i�/,�4P��2x U�`d�[�J�|���@�"uN��	�_�V]B�y ��C�	i��G'.hl�~%�Ĝ"��ˌף6����Aˡ�e�Z��K��_����{s�H98�`9�0˼�Q�m2E�QN3��@_M2��zV��02�'�|�p��������ŝ5�lu?�ѕ�a��������?���e_���Y���2�BS顭d�I�]y�Mqu�R-�B����G H�&G]�E��I���I����̀����RWH>���0�cYȋ�gz�f�宼V)�9�N��4����K�m�l�KWC���`�<��
�|�6��-&�A��?��c���Ty�Z��!����p���z��3GǉgIq�~�X�[�3g������]#1��f����ǝ;�~��^X�fO>��S`���3���'�= wF��4�k�ۗ�T�f�wpJX[����8�KA�@ ���"��/�^�;�f������~U�t�2(T�Pp�ؘF�2�Y�j�B�p����7��y�+g �>��)*�C隢��	��C�Q>Va+]�[!���c��o�˫���Q����/N�y�4VX��fӂF����������&GiV&�|�2�1j���$�T��-}��\����{J���䌐^�����؜[�S�"�<Q@�NY��/�&!{2s��{�A�v���b�h�ӊ�"��DOS1v�[�f7��7[�k�r�+�V�]���1��&y�Vh��O�|Á;��%(CG�׾]r��M�wc�P�-���}��K;�Gܓ����V��H��Ih�2�;v���z�^f&2P�δ1�F������3x��e�e �5ׯ��e?F��"�TT+𜖚\���u��
��v*k��2n�Snk��A(���i<��̩�P�a5�f?Gr�,۱�B�~�
��I�,�g��tքx$��i�{P�\��$�4�A���?���.�mN�ˉ��0���}:(��W�<��%��Z5�VނK���x��ɱ��{6LP�!B,Z�|;�8N�	GȂK��t 0{�8��K�Y�Tu�؊0SN� ���}�a����b�@�֕���p4ܘZ�d[��^l����c�z�,U_�7��t�+Z�~�WO�X�Q�,o5�/�`->��f�G��&�OA�
{FX������.�#!�KD;��b^�ߗ���7�%ʘ�p2L�_c$'5�U���ĕI�Ox�M�#�%�~��3��B�}�Z'�������Ҡ���H�$�;���B��*81} �柳�������zR NF?����CAUp��e���D�j�;>�ă�r�szفI�|?ey��!�z"ԍ;�~|W��]������T��Ν	Y+X0�P�� ���m��3�u���uY�o���za#�d�����+V
�ȧ��W��&UgR�"��Ѵ��>}�p��7�R���^���o\�{KW=A�����O��[�:�����a"�8�Qϰ�UQ�ZH(��XP%\�.�9����«n?LQ{�b� vyc'!,�(�&H���eE��o�)5�Ă��j�t�n��C�!EP�#�E�����l����;��i��1��4�w=Y+LQ`�I�4г+�}'7?[B���*!Ք�ӡӋ?��b�_"[�kl��*�蔼2\�O:E�[����Lr�(w.\V�j"eJDH��&�I�u��ָU��A�K��%��by>0돭��!��>�H�R�C�"D0����G��l�to�o�*�/�����vZ�gym8$+����>���Yɧ���9�il����l���0��%�*1Ep)��?����ҝ�r�ӊ�+�ܞ��4�$�" ����kc�}�q�E�+��>�Z��=�;n;c�=�YG�v�qϗlK��Z���/�H��74�v��c6
yǸ��H���=KA������7�w����>1ڤ��ڏ�f|��ʋ@49��y�}K�q�Pp�謁Κ<����\&	c�r�u���� 8��PT��q�aOg��N�x9�}h�z�D�4<Ojԩ��-Ф
o���:��K��_��d~�hG��5�AL)(@��YH5חVj��ڽ�v�����s4wje�8�"�w�4���,0=� \]q<�~:)��p�'�n�����4{+��Ⴋm2Q��ci`):XG�(Eu����#��G�{@��yN��l(��ЎRڥ*AyQa�PW����O����`��c5�W	����4�ڽ���Y�wO�����U-^v�Y>��/@����@y'�|C+��"�W� ����49�����]��^�ATauܑ���2��׺E�n�L?2t� mZI~���p�-U��*���@9�_���4�M���7@��3�s������H_/^m�������!�6����jd���\�p�eS�0�d>�Y�J�iY�#�{'�����=���l��V'u�9tؓc�z��'�0[{�*-&����>l�F餭s�&D��Ję �>Y^د$���Sc4?�d�J3��vO<O*�Q@L���"~s�o�t"3ټ��qĕ���EO�X5!��V�*�n?O��r�c:X�����>W�bw�{?DC�T���ׅ�[N���ǒ0���r�J�:�����|��⫊t�;jKp	o���P�/nQ=� �͉�͝(kк;(J�Q@0mq�;<�v_j��2��ސ<���V�JQ#z�H)���No$M{&V��B�`�wW^_/ ���q�cccb­����2o�Q�L=���j�_B|q�#�̢�a��R���༁9�h����ѻ�ϨE:��Ԃ ���^��]E)8��j�?�R��W���1`Ѽ�'��"ju��D��;�^'c�ʨYbj=e�����B�2���//�X��r�������G,o���S_���I"!	�	�Q)��\�]9�{-Is��Z�Yh�~ #�W}�f�6��@�q��4^ޡ���G�*�����D�__l!*Ҕ��AbObd�/�����MMA`>����˘�]�fԐ/�=���<ix�
�v�8��_@k�<Ї
�����O�'3����s��"�.9�ኽk�?E�qt��=�{�N5ɂ�J�O�ֆ�_I��z����E��f�!W�W+��?}��sk�݌a����H�䰹�i�)��&\�0���:�K_578B��e˨x�H(�*���">`9��ڑ��P���Ɨ�&hu��5�_ ���?�DOr�c
�������,���f�J��E�
��B���S������u�Y�j�?�5KL>�T�f�Q���_�:�㲐ti�{�T��~�x@�9(wU/+�V��(�T��+� �x���h'}�(ڑ�bF�Q�����x�J��e�QA,�q�A��X��n�y�c��6HJ���n�D�˅q��}�!�T�g��Uo�&��<6��`͑�l�\��`@l~����mL�9��Izߟ�#!�eĴ�Xѝu�|����V��^�^���=ʫ6���`������oA��i~w��m�zG�;Ϡb�#ZK�c�F���Q�S&�'��-���ə�$(�;��HF�GO<��>���4?�7CL.;�]:C(����	#%���$Lo�X��Qu�� g����iT���{k=���������va�+�y����-[1�0B�����t�_|�\�È��՜�|�2�%?�z0��]�ڭ�t�t���XɄb����p<�������nu�w[: ]��0~e�F�c��v�.o+��b�H7�6��*�B[�G ��Z��&��y&>r�˓��	2���1���$v��s�����<P���<��j��o}]��~�0}�-	�!��: �ӫ�m�M�ך�m�!wǑ����+�Zi{��X;�^��6��+{�s� ���/T��Y7��{����?W�my#@2*yS��T(����5���2��+`��� GN��}�s� ?1��G�j�I��W�������*o6����,�9M�0�қ��{h��ʌ"��c�	.� �x"�у�ox�����,)�tCNRT��5�Q��N�b�ڃw�B�o2�B~<�n�����������%��8zwe�'��  �:���A[��AߨU�i^ܣ�M�5� �e��
��(�\Pl9��*>;R�Nu]Z� �N�m9���}ko���*z�\�;�[��ve���?����Y��C��4aX��� w�b^C�p�
��g7]Z$ѯK���~���k�����rU�Ҏ�DT�3ӎ�l������{��\�O�eǢIۀ��,���ҕ���x����D/����rģ(���zxY���Gg h��M��7��XR��6�/��O�SZ�.�F��]<��"�4�[W�p���>����^[�w:��I��Z�P��e~+��f^���ί��2]�r�)���[3�D-�F�w*@F9yM:���q�"^����(�%�L��1��X+���Z�Y���75��zjtD��b8� ���tHA�C5�|�8����ʂgN���7��ȾAHSujW�5�����?]��shaNS
g��R>:	� �`��J�U�3ie4�6��p��"��Fbk9%��\3�Y?�������9#A�|fg��!�Ur�5�͇Q�/�i���^�o�͘=F*��`0�v��h�o��̗�(�V�� ΞRR�4��X=a��e�oP��/pF
�寫�Ǎ���փ��?��%1:����%6oO���
��B"ca��t}z� B�>�R��+B�k�!ꐨ ?�u�\6�A�����c��h;�� �3���B�#z ��N|å��		�d�P��dK+A.^�x�����Vt��q<�+���3��Ϧ��iH�;o�Y�V����D��%�e<5|�j��� ~��{O�S.>��`	0���鬩@�g��r3����Ն#=�>��|Wi���b��@F�6�rHF~T�UP�ϐ=��[�F:�b��/�w|�2�s��������Ź�V�ԃo�jh���x��#��#�})
�k�n�É������y�X�g�|.�.U�/����AUS�'�=}yGjo���F{�����
�7��EQ8�Ȑ��ΖN'<�"S�4����Z5.���w�~�@blq�)�qd$X)ו���P�g鈳
�1����M��if������/�kU�@�ʐi?a�¨-�a���W�@z+��O86�ɩ�r���a�dp�%�[�/��o�{nx~�}���!?�\�|�[� >S���|8a�S�� �)�R���C�!��:f�*mM�}���r~��Ce��b����0�sԠt,L���+��9�= kl
5)e�F�ƺN��=��� ��N~�O��@�;��M�>��s3��C�a��*��}����w��\YZ\�\vRʔ�k�v���G�<�F����@��X�uC���tBnJ�0M�����J�o[!7�_���GKg~Hf�@q���=^�̽4箢��K���&����*IhR�=9��R��̶�O!���(�B��u-7E�[ ݡ�>�|�&6ς#$���/8���<�x���L��N@��PE�����a��-�a0�����ؒ�T�Zfûi6O��#�?��7��~c�%��a�K���-}/��脂ːH?�e��qw��+ۭ��*����m
�8mPWR�;��v�~ ׺�p���{lk3C�HH��CE��̚�6���KE\yZu�o���_%���.�[��q�����^�ʾ�e~!:�g�ԁ������,[����-��h\�fFĖ�;0�A�)X�31c�u�D'���)c�1/��MݲQ�㥂�9�^� #-(�J��@;q�����ǔ�Hߋׁ�^F��7H����dzڀ;���/���Up1��C/i�q�a>I����P߫�fD�d� ��w�c�VYH�t���2�����e.���%�,�+(��������5ݞ`��S��"α������Wu�C�Q��Ty)tM8�`�� Rϼ�9��Gf�@�R∠@�c;� ǥ�Vgn���/~]����^�������T;�@������KkM
��,�f�Y�q�c�����?;
��7� �镘�+�v�x����(��l�C��}��7\d�ZA��B��%I�0bd�&����1���a���]ǋ���1�]�^+��!)t�}��Mt�'���U�wG��F���C�=
��{�	�w��0d#ѐ^Œ���c��@�����DV��/��y���n$Q�5�En��E
�|�17#Y�+rn�C�f0j6�˘�����ۂ��I N;�pq�~�|@h���sd�k�����1��� ��*ϿЯ����,�a��*��J��
�D��j��q�:9ɕ��b_^���Wq���%��?���n��:�8fP_�����df��B�F TN)�d/C-:cD:�y��kf`R۸&V�S���?��E��@Ȳ�� ��������H0e�)J���uiL�c\ܛ8r�^I[A ,�z4�C���ͭ��rB��CT������oˀ��xBj\��^��`$:�ݽ��­�fq���/��=J@���O�?۳��HI��?��#D?Fe���������]q�P<͏O������R�2F$|�!�šD�b{`�fVqL<
��v9u;�.���8�$��o��˥�eY��qe�\?�^�B5f�s�$OE`9��L�f.:v����2/9�,w{UA��2������-�����=D���բ�u�a���0�2����1a��?3��$��k�W͑w��P7��?���0�_�E��Ų
=
K
B&/�f��v-�'��	�8�6!?�>�&_>�A�4Jl���3�C��6��_���QNܬ�s>� 
RY@=2�>И����'��pD����J����� ��4ګOf�@Y�������"��#*��Z/0bH������Y`R���0���I��
;EC����~�4�Hn���MPa��:XQ�P���c	���Aq���5��\�{�T|��t�i&;-|��&��|���i�������d�|��sF�g_�����X��x�z�zӗ��<�f��ng��D��<7�E��]<�6Ů[+8�-i8����S�&�g�F/����(������7��a5�@t����2Y���L�` d�g�Fs���C� r�eѐJQ�
�����������	��0ZP��~��Uܱ�W��[�$z�\�����P���B��Ui�r+A��Q�z��\������g[��U�<Wg�?6 �Wֶ�z#J��T �<���~���LLk�m���
���7k@�)�ꅴ���\���YY7��j�g?�D��,ü$�^�iHP�p���Z�i����)u��,ƍ��m��n����Zv`9b�vI�+ƕy8"v��y�Ŝ����=���xi�6dTX��i�$3����*F�+:/�}��K�A*�n�����h]�R"�m��+(�f@j<�����/7)�WȇK�J���SS�Ӎx���R�֝�����rF�)�1�/�k(E"c��-���oA��4���u�nG��}�S�|�f�W'�A�=��dh�K���t���*U�ђ�c�5�����YFݼ�W������M���� m7[��������\.���}��Őu�U��$!($F��U8�h0��}llv�a�K�Tˇ������7����N�:X#~�x���N ��*(�_����n(�d��'������,�X��2��	FV-\ǱyA���o��[���̒�#�5��WSb�dUA�r�^���xc:-s����.j&/�+�B�̰�z-�\B��L ��#/$V�-ļ�� z�����$�ǆ?��gfs��M��iR�(ypmfv�Fo�~?��pWH^ ��ƇS~�*���,Z�/��t�+x{��i��K`Y��U~�_�h��!4�Y��]��ϱs�H��_a	��e�_��:�>�גY��a�Xq
�����\B�w���<��`��Pbo}�'�2 ���1O�D"p1�Bǌ>]�B�F^������&��g�gVу��=��`X���1K�3�{X1���s��ß J��'��U�׋8N䢘�V�$;1�l�^gUG�<��ݔKI����<�[�:��i�A����!zQdn�8�:,�Zk9������N�<�$�Q�(>K���))`����R���]�Rjgx~�qiƉ��6y��&�k��lE�44"�.�a���'X�.�z������Т2C��鱮�_���́"Jw���[�_��7�}ĳ6��&e�2z%�W=ݏ�W9BQ���68$]�M~�!j�l}ɥ�k�4��*�@(ļ%�*]���J��Y�x,y�_B��1��I�Mqs���:b9�D�G���L���b��F^��B~�������n��f��u�3�5U�ܭ$������\m�`$���i��]AhUb�wc}��k�%Ͻ�!�Eg�R��\e�`�?����	<Ph�X�̗�\��ut�"���'�U�+t��	 0�b��Y���;����P�Ţq-��LlYY��
L�I4-f���T�Bh&��9z��n}� �Q~)�2�fS�*�P�����g��!p���l��O�[.'�)��� 8���e�\�1�����k� !P���M8��e:��$?�d��ȭ�{_$�x�q�5��͓Ւ-m㕆�����O�lPٓ���&�U3W��� "Mr�Q�IC���%� ,{�������,[B]����l�KX����bX$F
V��G���+���g)��g��,"�Dm�}�V���T� �kF�[�9��b�,}gG���L.qǏ��	���qE{��	�����L�����\.�8�ނ�Q�g���UT�|	x�e@�lR�/~�5��s<y o�2S	�?�2�1�S7t#H��1mq���z��Y����E&�b�� �)�

^v�HvTI�j��%���嗗�d-P�~�ͤm\��=�`���P�c��+x�uG�KxC&TZ��**��?	h���y�|�����A.�}\8?H�FJ�(�;���F�I��|�f��h���?(o����W�G��5������j�iG���]axT��ze�F�?��7Ă�)v���$��k�+H�=�C[{+ﱷ��`�kPנ̘ypJ�>��b�cwqh�vHj��Q̈́��NO�톬��Je!Jٳ�A�>���v�[��yt�NKXM*fű]��S]ʩ�}c����mw;b�y�Η��O�&C�ۧ�Q{���D�sB�}��E�|r���
��A���ں$h9�zu+������@�DqW��o��o��Tg���U��]��]Mڨ���hm��g�a_Vӿ_�oό�%i�	Dk���P������uOa�m7r@�YI��3 ��"��L�4L��D��@le�KT��KN ��CުSi����\I�U-���}=M�\}m�d��y������8z	=P%s��>6}������B�'O&�T��X>W��� ������$�VGF0�"V6�?⍞^J.�z�~�rkf��-yB߼�Є��3��FtIM��Bz5F����60_a�u3)ޒX��ޡ����Q!�mb᝶gy�`eD+���~[@O���^m5Vi������;Ab)�L�,��l��Et恣���8��p�y�-T�t�ϴ�Vw!2�Rצ�Lۆ��PT��y0�V:j��"@���Z��|� ���bP#(s�)P?��ӓ�v��G5tyZ�`�aG\,E�Pg�����|ua'H6�A�^��q:v�ʪ���OTq	�S�3��IF�Ș��q�;�N����gA� ������op�r3e�ټd�ٶ΢f"̦���i�\�Ɩ�՞���EmZq�S�����=�rc���:z�:(�,i�3�X`�2V�D��g�ya&�7㠻5�VەyZ~�0����1ԡ j��.���ݺ}_�sҁ� �}�?�$`�� ���F$�S:nrs��ul�F���|D�RQnL�~�x���\6 ���ȩ�u�HA�:ģl�P<�c��|�%3�2٢���
��r������<ם��j�a:��Ћ �q�GkUk�(��߁L�^8&I�/�92ն�ҳ*Dd���UF�E,�9����Q���5yNd�����ag�«m�Q3ك!|������;	e^��)S��?��1�`+*C���b�o���7��GM.��k�> {�'�yk��z�$N&���m�%EI��%�s��E�4��*���N�u|y��(�E�s�y�rݗ��En�bٻ�2#�����rꆉ"�
A���]�n^����_O>�`ȁ���$L��x��?azeBc�66��Rˣ[j7t��BP��䥟S��\2!�y �Ȯ)����鵼��B�+O\���@A$7QS!�A߳��<n��J��o*�*�8a�[��`�բ��൳�8��TW����V�
��~�Y0�1
�����Y�7<%[L��#�k-u�*Hl���k��.9�����
�N��E��'��Tw�K0��%fQ��'@��H�VO�y�5=�B�A�B������Al^�$?���0 cꌺ��'&q��w:e�*�
Yi?�R�C/�f������x���������F޽xe;��e��g�(cI!
�����1��Ԓ�+0�S�oWv���IQ�\S�c �[�-�a� \u睙,���ܐ���5��t�"��8�P��!�/��rЯ�+�$�Ŧ�L���1�j�m�0p�&�Rl[%�G2:�ǋ�.z�I��66렞Md�2�FN*���+�縛��cuݙ���T\3Ul��E �х�
b���Z�
��8�`���C���ͣ��1�a_+� }�'�ۛ���7Q���C���E������d�e)4jh%ë9]��EV��8*1]$o7m���Q0A_8������נ
�U�.:
���u�u37�@�����
w���NO��̯�,q�u�J�2���+��ԺP)0+^��8��Hp�TlJY�w�]��t��/�[��f���R=?�w���1�Y�_԰8;�k���ѱ��<OG��1�����Ҹv]�.��]��"|��ڳ+����(�6�
#�A� hR�� G8"���Ӿ2+��S���b��"Ԫ]�����|<�wh���	#ἄkO����-���s2qtRS��Ms^Uf���I����F��ϓ}78+�"�J������&��YN�W�r�17����{�vI6�'6���)�x2$;�	���m�T	@1O��^:<� �:` ���	�z
�)2��E��?<�~ɠ�l�-��h��?�Ժ�\������̖�@]�EC�y8��d��+�ܖEH��9�b�}����6��hq�o�V��R����3�h�J<��ѪE���_ ؒl�M���f�y�Ps�)f	����M�뵕�XIă�^��(/����j&1�zJ�Xx�b�_��E#�L�:>��{�ID^p�ʻ���i�Ⓐ$�����fǋ�3�4��A�	�zrc-B:���j��h	j�>&h����<�LZ����`�d\���H�%ΦrGۼ.Y���n��!�K[9 �h��h��O ;��lL����U�9��I��ܫA�� ,���Aߛ����s̱	n>ziu\\���e��>/��ȇ�����VY�faB��_L���n���I��-h�7�����͘Ѯ=妄��M�M}84 L�	���RY -�
���� K�8��	2fRS�AM��t�S!+܅�7	��_y�ʸ
�w��.v�k^�%�G+�ѝ4B�BY�Uv�їδR�'z��V�u�H�ک,�>�	Od��%�~q��.0
��1���|_��:?��G����ܬy(�Z��f�'x�ln�ȡ,nFd�sD�P���Ȕ�����e�Zv��&��S�iy���Q4|;�D���]�P)w����,W�I�Հ��[U^uFӶ����~Ki����<�B��۴��������7xT;�@�:5�5��]�>&E�����vj9�^2��6�� ��<p�'�T�w�$�PG�X��{:��-՞�����\#��'���ֽ�
@�6�##�p6�&U���&2�3�ͪ�)N��k��c<�l�xT��5�e�*��/���F0IDx9&���Va; U�V�D|��MR�U%vȅ(P�ے�p�+\��곙�0l��ۀZG"�U����'�1��+LU�����!��,��M���)�,|�����鱗ͱ�J(���	s��w�+��f(����^ҫ�ߡ��N�k�>�ZqUտF���|'�= }\*��}OV����{���$��$��F�,K�1�Moq�$��ꤥo�p�Ώ��X���(t"�X�gH��;Z�x.�˂�� �'�*$5.��
��t�G�Bo�Z��v�u�2�~��Ԧ�[�e�
7ruy�^ӨT�$��s���=RREw6�I=��ؼ��_��`��}E��8i�:�}]����tf��k��2�|�õ�pPy��7�^�J� e���4�ſ�	�M�kx�:�� [g���������l
�Q� ����u�E�SZVT��Swa�C�).�Y݉nh|���b��mD�Oޑ��ǻ�r�|P )�4(�BF5^�цpsm׎{���2/�̜0JԊ^���5�x�$�?::By�������Xd鋊xM�w��?��8�a��z6j�	�w�Lnޕ�#��o1�@N�-N�="�G�K��gH�A�<�=�私����TK��)�V������������گd���:Lr{A�a
&���~��[)�%��*��n��� }8��x=Cτ�3:�Кh�
�D#�sL�ꃅ�W�s��l:-x�Q&�����
Sf���8����i���?�q]���GsgXNb��׀�hsC2iN��q�vw�?���݈}j�ۑEk�%��+�B<�(}u&���\z9�~���e���2
����5��d�`�bс���v�������h�a�[�Ź�S�,��=�V��F�+�AG�x@\Wf�Ӑ�����4J�j���?��9��������T�;�{�(~��H�Y#a%KvW5� Wm�#V(��_IQ?o�U{�?���0��ז�d3�kQ4Tb�s�p-j��tY8��3I�)M�7?��?���:���)4/�j�iZ�P;X M�FZ��w����(H��55TCX�D��R����<H5��U#$f�z���9=��`r�-d
6�ZB����K�4�'Y�R�cu�~*���`b�b�;�l3cB�f���|g��:mhW5�ۄ��ggŃƕX� ��2�s�@���h�#��H1�m�@�����/$��%4}�4c����K�� T �����O��F�9�aå����8��Hv���XX�ӿ���y���9kĊ+����:��i�s��mg
��&�:��)��t�CxU]��!."#aEH3v����㾹n"�묭՞5N��@Gat��橲%�t�F]c�Ě�9@FZG�)g&֨���ǟB=�:�C����-�U�p��J7/9����`�-��!my��:U��� �@��Q���0bc+̪5̱�=8p�}&�B�tx����c@-Z�*E��H��;�x|'�Y	C�M�-�]�h�U��8ol��wM �p����!�����\}�[=l��bیL�ğ��� �慸I�[��`"OeX�'A�,�iE���k:�X�g{vƃh>�~�XQ�D�^��R����:���ݵ:H9]�º�rSl�|�`���S?�18\����Y�gUy��B�i5���'ŋRq�qbo�~)���n�g�f���-�hy:<}?�?��Ή�}�Aܿ#6
^���<�K�66�S�)�C�����h��n��E�TB&��M⠒��30�ũ���o�[3KI�q�����Xa�Ӳ0�>] @��1�i�";���;�b���3�&�FI��m:�Ģ�Ggq(���4�
�M>��	Fl�a�\�c�o���ߝ@��Wwg�ؓ�2� ��zo3��To=��u�
�%��o��y�p&�\��QI����,�b�,ֆ@x���6[�#�@��� Pʈ�f�[�^g����B�/������傰4�GC_'�>���B���Ǖ�:�c��c�D�6L��j;�C@�7�A[vdz�AvY��u��ik��7Q����:?��]e�����Yh"|�T�Ѿ���n�����ϋ�p~m�6�z�
�	����W�_e|��������S�M �Ղ���ic�w�N�)iaFr�����s��aQ��}�yZ!�~��ꌔ�X2�ځTr�w>2��%�Q�P:�<�����&�H���j*���AKqX�Q��e�޴��6/�I�*h�X��ʄ��aw"�{ ����X�3G�Nr�O?�(\�G)!4#��wNl���D�$��u�d(Wv�j?��qSC��V˾(!(=Mk�[�4u�V�*�S\�<�]��O�]�BF���,�^�;u��1q�V)�8���=䔫�u�a����@�&��11aF�Ԙ��F����Q�0D����b�'��j�QNv�<��%0�{��A�ؖ?$L���{<6��*�	)��R$��JS���=�d,ć��q�&��L ن�Q[[c7T�<���4;kʨOW�PB6@�+"ff�ni�V�T*"�{h=��S��Td,����})ݪB�CZ�L�7j��>�\-$��J}sq��c��rd�� %���T�1��� �Ah�^E��v{��L6ӿ�3Z�b���k���H�7�l��l�+��ė�'N�!r;r��K'&��yQ7R��҂.>�&��u_��n ��md������ɖ+vY}B�7�>��<���Ձ�������� @
�ߔ3)B��{��L�"Ǣ4$k�p���#
�&Zuj�G�8-v[�Ϙ���n��d@�<��y�G��L6E?;�7�:�Y�0�m���`����C��ez1�8���1��Y��aT�̷�Y��Z�����m���t�#�y���Y"o矡��d���շj�����j��)��I!������>��S	'٩(N���Z�����u"	R!�>�[�`@��ȅ���J�2M���@�����"�E٫�A��t�MlA�fkl�����B�L��6��5���W�^Mk�֚z�=�ȼć2It�H���$��}���i	��@�����5ͭ�'�ݿ��ZC��&H+,宗�:J���"P|��q��ZŐ q6>���E&� /������~�QR����F+=̊e.T�GF0��
gA�s�\�"�U�����d����']�`Hր��+4W�tzJf؞N&Yȑ�0��G���*��6oω�g�w�؋3���-�2��?�a�pyf{�,�wx0�?N_*)�6�쳪y� ��76��s*�#��6X��N���y�ƞfFV�E���+{^n�opXe�O?Ș��A��uc�z���Sv¨�/�����\��� >/�5¥SvN�{�1��d\�� c1���O
��F)]>���sC#�a�0��ꕙ)Ey��li'-ɽ�����13"ݰh�,�"�/��R��8@2íS�[�'���w��";E~J�#�~�J���>�P1�Z��Ҫ碚1��<�L��ZW'BZ�!6�O1�P�5���&Fה�*�>{�>�o���~��c �^��+4 ���9v�s'���a՛rU�3���~��e��H|O9U�t�o�%�k���´o�jK Hz�H*�����z�X�E��OSs�����ӧ�̵��V��3 �?��xp�VUc|���f�#rf���?����l��-q���2��F�� �֘|խ
���ϰ���P����v6��
���p���B�0Z�T4�%*�q�\�{Ǜj�&O���}�N��گ4޹1._^i&�9�<��~�1o�����A`N�/����$�s��<�m���` �B�\�!\���>�3�05U`eL��ݲ����3�e0��BMRtX��Ie�=gIk+kr��x����� �S��ڬ�h��Ճ��[x�<x��	4�逗5 f���۾nr�+�~��V�H�zĵg�X�P �����ƽ-y�4k4�J55D��I�x�hZƵ�։�������-�^=U��og��x�u9*l3q�&�dPM	!�'݊�i�H1� ����a����?3ͬ{���Xs
]K�j�an�� .,;���:f��(4��x�^�O�Q|Y����(���p�R��;H�I���K`T�߳N��V�,@:�N���ӈF$D�3�I�������78��cU�0OIT��o�x�R��䧓�F�G U�2�ݴE|�*J��k�-�qלx�z����U��66%�=rW�+Y���nJmN��(r=T���F��CP02R+�{u����cgt�P2���w۴���b�UѸ ��{��&�U<�����X/Q܉����l���}I�p��;�YU�����D���Lp�����H���|��\���Z˯�ǆo_|>W�'7�k�����!;hiu�/���~N�C���Xh��%��m���T6a5Oj1�/	}q�Nl%jHZz#O	B�Ѥ*[IlJf5|��J6�Y"���e�5��xƷ��*$�b���J ���z��QQ\��A�>,�9��P�S�'za�_�j=�a4��y-��0���m�8ר4���ud�?_b�~#c��2�L��|��y[1�>�Ř+^���?N4b$�YXs�^��#��
���)�C�G�܍m��$L��-��s��k��sSQJ��0g����s%�.}�P���'l�3Yړr�|�]�p���Jόv]W�7�����8�L�umP$�&�vU�F�W�>o��E\-6���N�qѼ`�h���/������c�}~f�E=,�-!s���� ��W�Z$8��b+|��O1c�v��D]�D�.�� ��/CY��sQ��Ϭ�������2Gn�W�Kn�a����Q���I����W��D5��!���Z��_<�����Z-@^3�[n�]y!���2"�BK���rOj�{�6��g�q}V��̎t�ߢ���)��D;��Qm��He���*��4M��n�?�Q\��<1#�5
