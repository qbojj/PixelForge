��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s������`\�3�*ME��!M��5qN�H��,��?�#ߟ��d���&���n��
���XiV��	r�� �-|i8���vꬎ�3q�yپ�;lV���|Մ�[���N�~�*�yTL{��+Y�4������7Ƞ�i�ޱq%�VW���B�E_	���6����;6�?���N�>WQ���x�q>��a%2��uV�O��
�r|���Gٙ���Y�Â"$+��:�>��v���l�g����s��:�h,�����Ƿg!�O�}�n�$��$mj��%��%$���ۙ�mܓz�,<)ې�+U���)עvoT�� ��V̲M��b7z�lɰ"T��hg�����k����kԜg�9{7���*|��W�`F�0�Q�����}O��W���ZBj�ML�P���;�b��ƈU�b�}x�Q{~���D(�]��ۣ��_�"� t��#�2���e�K��(�p�2'ko���/P=pw�a���!Tt��W�PU5[�u╯��EE��k/�Y�
�S��P�j���x�,�)��đ��)�[|k��߂��|�-����e�i�Z�<�� )Y�,����07�F�Zp�\MI�(��故][Y��3�d��w�
I��g��9 ���
^l�Z&a ��д��"�=DEOO���o��b�l�/>���P��o���)IR豃��h3�q���+㨋e��Z��8k!�;iJ7Kg��n�f�j�z������ϴ����˱�G�/Z�%���8�O����~�S]�1f��!}���J�C���?#T��JA�}4Ҳk���������:��o.��M)��q/��LG�̨\i�H��Y�2_㿔�tȞ����b�����P ��:������X�M&�@~r��~��#���BW��Џe-~]��&"��ak�?F,G��/��y�7\��'p"�����V��-Q�e��.۴Q�/�S�'�>��i�/+��]h�#-�}��L܋s���۰�$�b�+7�FJ���UNqERսz+UƚM�b�<�\?��9>$�"��79��3du����� �h�N�����ٹ?���&��Y�� ?���g��pM��y��u�/�R04�aN�}_.GčʃB3�c��U�=[�(��-��1�H+��+�OY�h\,IX���9ߑ���:�h����h��ec��#�9]/�]����w7W�KB���\ئA#c-:�3'�/+:9�� b�É��(�#}V��s�"�$�7�g���@�x
(��|pǐj/�:��x�';+h2�(^D��gC"$@�1x(��w�p��L+�t��ݸ$��0���Xr�Vv�������.����f%im�ػƿ�t���t�eN�ـ[��}���ɮ<�`>\��)1*�ʦ�B"S��J���6A���tSN������ �O�w��vBt�s����z`!�.�~ِE���h����PS��%ܼD�	q�C��5K^��|kF�Y�۝�}XI{�_��#�AЗ?��xUw~��;~�Xh��/ŗ�yv��9��-���9Rp�)��M��.��H��3��+�_`uJF]�RA�ZE(�����a�7��7eE�c���˝�GD��S4Al*t� �ꄫ��O�:���8C�>t�k2�������h9�it�]�SŹ6�b�SAL�܋qG�i*�P�^�6��$t�dC���I���[GB��?ށ'�d�f�ݱ�:�Q	fъeXĭ܏٬�0��Kv����fqs�?:n	��y�qѸ� �{���Q)�?Ś���6�k����(�a�DL4K��؛�rﺂ�}��t� �b޺Ծ�jl$���'Y�b!���p����,1�r�y%t8���6��ܝ>3t����H�̑�
Ƨ�a��΋���B'.�`�N�Mc?�Rz�6PBb�ہ�[tq�X(�#+5�oy�Ij��JV��6?6�2�r��"��%#�5�x<��2�V;�?���ɴ	a�����+�n�yW��H�Nfo�}&��q�'L��uR����ܻ�^�qCF}*P��o�U��Q+���z�	r[4�!x�d�ld��~A�8aoK���X�"����W�ւ }�X�N���0�s"�t���$T�A����e9�N#\Y+��J=�P����e'�d��FKLd�XǼ]���ٲ�<��� ��߉����i� ��i�$�){O����l��uLS��Rg4�|@��I��eS��8ƃ�ڻtY�	P2c�[Sz'��e��[W�\B�:T4�`�b��3olN<[M�e�������Wt��)i�E�ΗJj݆�F/̕�;p��.�I@����9�����&��[��+��ɔ�N�7��:<���տ �wY77Yݿ6�}�H1����<�������Y�e���=����k[F�t<����x6|���f(�<R���J>Mؤ��xPO�W�H�H�K��*�e.�`�
�ؚag����
|!�18�Î$��3Q�� ^t[H�ۛyy��-����>xi�@�6�V�)%OJ?���H}��u���/����Q}��*�� �[�5V$+��]T~ߨ֭�lAK�}e�[���v���Q�}���#����#�}BO��<>�VS��pg>��ǢL�4(�?_Pf���� a��jHy&�M����BR'�� ۧ8�NIj�|x�xb
/̪=i�#ϊ �:Ͼp�e�k�Ƚ�&H$�c���]�|"�i~̛�J
AkFI����N<�B��m�}�C�\0�يɝ����2�=PZ����5�a��A�+ў]+�t��K��aqx&g9ź�>�+�2M�f�����}2��#���k;��j�+�@l���#���|>�#�f>BA�"ܗ�)=��ŵ��lH^�m�#���T���"M'�W�
�~�O�N\�����Q��0�U�֬�lL�9�i���j��E��U T�!�~�{
�����w	!�u�J¸D00-�	�	���֏%(��+%l�W�B�t�έ�㝂�
l��z�p� }H@�c������f�k�p���|ie�O(ǣk�u=1�gS�2��n�?��O�@�~��[փ����F�1���!��Ѱ٘�$��6a���z�Yg/8UY��د��B� �S��raV]]�m�!��4�q���~ C���5���L��F��F���6��^������Ԋ�>�������u�������y@u�N�ZV�"$��c�7�im�?EH{1$�v���슸h�K*�
{��Z���i��kxVc�RK���=V��l�J2�9)7����b9�9f�"q�!��-I6C_١�a��B���W{-pAA�/���C�|�B7��Ycg��WW(���W�Y�Los8+Y] ;Bk���]e�{������V
��w�?�N'"��G���x�?N�����J
��h%\z����-vOcٺ�d�I��7"�D��*�*���:����>Q5�W+(a�JcW��]*�9o��J�:�8�.�Tn�8��qE��0t��1��e�@y�r7����������-	�r���oH��b��I�8p�	�C2����2(���K/��ϫih��Ef	CA�@��8�[��r��/���]d��-� 3,���!�q�U�;m��%!�Ĩ�oש�S�iY?ݯP/�(C�N���]��:_�*�%�ũ�mܩ��O��.�[�l?
1�������h�E�Ϻ��\��PC1O��}�!ti����#�����\�jQIj�(��6�%�Ǽ�J�#���]��l�	f��h1� ��杺@������78#~G�)c������W�(_+���7�0�z�?�X�����ݮ�H�{X��~�9�/O�_����~�Z�[u�^�	�2$H�2�B_��)���$�ge����4��a���{<�U�y�B��q� �4]��-�,���Szp� k��%}�})�hP6o�l*�ea�~G�vpA�x�X�_��k�M���X��ъ@���WuƠӟo�(E�3zJ����X]�r��w֣9`k[ʉp�G�U�xm�Ñ,��-^=���#>��[/�ٽjȷ���K�}��$"VR�q|�,�9"�|���Q�Ф��Nt	�<bl���c�$� �����7�Ű"���gj ��Tj���T>�\�ǰ��?�ͤ�M9��fxLP�����8U��D���NilD�bމ��o���0����P�
�Kk.˪^�4i�;�귝V�5d�`����
rl��A���3\O�9���c\~HT�R���O�B���3U�]�&J��'�Tt��Bz��^ğ˒ Y��'�Qr��-�Uvr��U� FH��2%����s�䞟���Ts�0��R7�ߑr�E-v�cW���sv���
u�SyYM�C��E���<��0��i�9=&�����R-c3��Ś��W��<Y]��%n6�gJ��k��m�}�$���!��b�s���<�gHNTM����L3D#7�Qs8�7�[������Aݤ�m��5��7��`'���t��=+�J��lL.&��p��bC$��:���6Aa�A���@����C�����?��vʒ�b��3�:!�l�7E"���Kf�s��yV��	`y���|�?G��Ov{rB��g&t2o������W��j��y�.Ʋ�jF �_����1s��"�Q)�����4����Zς5��fTD`��Qr�$!��@���R x��!�����4�`�2��iVyvi��ʪև�r�$cR=�R�a�O5L܇⑾��Ϻ��b��!Q�G�~�!��F&�;�]RĤ�d#�b;O*wl��*t�=[�o|�0��A��z��8�`2 ))ز�H����0Db!�����w�!��c_g%P�팻w�5
���� |c:u�oN������+Ne�_��ف~���q�E�SҎ�j��r���ò�d�0n.;���~`7�<4ʰ�/1V�ef����MXqE�o�ꩮ��B�4������e��Xˁ%�c;�tq�4bC4c/��?7�d�aܟ47��_�	;�K��M�N��Q����m���v��$����O�U�Ve!d*+��j�jH�oԻZ�iЂ[�.lU��3́�B�7�)#R�8]�����\�h!,�]Ϲ���X&��y��dsT�]�j�~v��hc��*���iUѤ�<�_�t�!��mIt���x��H��`@�MU��s�"�9U���ȲD$������~ls2���x܃��R+�8�z���F�%��HH7qE\��R*�AS �'>����!�w9�-��������0�tw+����u�H��1�-��:������n sC{�U�ZW}� �!B�DlhRȫj�H��h`��*D��톍Msb�&�K��1|ȑ��J5��q��2��yEE�� ��������Ǘ�		|cF����K[s�E��8�X}CSMZtס�#�tld�yD"�4��?����?t�G��N%�ݐ��ŗb���l�S�.J+����
U`=�NS|�:��:$n͢�����jCUQ���y�w�-���e�%�Ӏ�L;��<��Ӷ��q*�j�762^Fr�a�K^D�x>�9#��R�$�FРKqk��{UZV)&"��CsXb8g�1������v�6`���p��/��X3���~E��)ަ��ڛ�*����HeiP!x$st���M��*Е���}�P���.$��"��-���%�3rd����6^o�Ƴ����_ze�M����%���IG����l�����]�eW�����AO�\��'ߒt�`��Ut3�/v�� ~��a'��ׄ����d��q�)8� q!1��:0���e�v�'��i��-�{n��L6m1����Y������j��T������Cxܻu��XXƜ�c�WÉ4��r��{��� E�B������[^�l+�{��f����fs�G�E"�>�H�:|�w'�����H�F���I�V��tҲ*����&�5���� �!Y�� 7z�<��MiQM�$�A�8��ʏC�}/b��������T9M;+�Z-%7FG�i3�Ez'�G��!aC�8������g�Y!�޹�`�s�K	��!ZΏ�	f��@w�B��[^t|��U��"���J���S�O���,N�t
���b(�x)h��,&�K��a"7y.&b{5�e1��q��s!��E������p��N�E}��f���V�����/�Q��[T}����7�J���0�i���~UnW�/ϫ�S����f�y$7�gy#7j��Wx�w�.b)�"��H�w��F�R	��'�����g����qv��G�D�@ն�p!����<��Uj�*�=8�s` "Ҿ�6�Ы8�^;��kn���Z������QW!�i9����س�������"�8�T6ٻ���Ρ����k[�B�j�*9�ɇ���IoVj�>�R��9��툩t�?�B��~�-i �L�p2r֚�`yf+Yw��p���$:i��M������͑���x.�^��w�f-���8g�XRȺB�'.�\߰~�zZ�����*Y��S�#�|u�HQ��,���Yn�I�l����'z��/�/�� 6X)+<��kC36��è�3�+��n�Up�~��H��)��Fw<����@xO��2vi1�>@�� ��W�CiH��9�� #4���dq�bkK���:���"�˚�~l�g�>[Z�\�nX�UD�6lC��Dlͦ��I��v �!,�Ȣr���z�z;�gٟ�bS��1��� ���j�+w���N�_�m#��7��i�����]0�8帋��n[PyKT})�L��*��l�E�lc:�A�p>{��tk�n-�d��c)@��t�d��mY�PR>l�̃�I�'������z��诨���yl?�e�ߴu�rm�NEY�+�`"�[�3��*P>��e��zQ��=%��|��Mmm7i|��L�
�iЧE���=7�8�I��"TJ��E��7�������av��|QQy{�F��ߘ�R�E����*��Ҧ�eK�1\fb�O־>1��?�K��+˙ٵ��_)�p����x/����PYN����RKf�iėa�� �E2�~���3x=IOX�y[CG�t�I{��q���n��M�u�沼2s���KS^:]�7�X9��tW����y�n>h�n�2�\�:���߀;e ��NA�u�"��0l7>�Lod�wm�Ϩ�V�u̓�F��{�߂ ��+�ԋ@�٠���a�k�u�N="K/�y�]M�7-d޸�`���k��eeNsJ���-#A|^��
g U�<�O������ �,��w��٤b�SUŲτ�F!7g����T�*:0���Zn<=QQ��c�Y�j!Ԫ�|n词��r�i��J���̔6��M�G���m.���=X��8$Y�f_��١I�a�>��J| �u0А}Z�OL��ӫ1O�L��n"k�C�$��s����,Cx�<�n�w�A0S���V;�C+]�,쵟ĩr��)�$k�D�O�`�|\D��&;ݬ$��ϋ|��j���o���s�eS�/���%�)@d�A�EcP�w��������V
A�z��|��[��{�\�����s�/2^-B	��Wycty������ػ݀��f�����m���<B!>�)%����(� cD�C�^���N?*���?ڤ�.�����ҵ�W�0F]�K�fI6|m��`�)&$@Q(��+1� �k3�{�{��4��m�T9�Ɍ���/�Ox3f�1�V��L���b%ά��&*a�"�a"�5mŊ
I�܇ħ������.���{x�!�eL��"�1������a1���.Ry�T��k�QI�\*��7]wk�?Soj�n��ɝ�ǈ��Ӥa�Q�mPOC��)�!��*Wƴ�z,gǽh�������A4�i�b!����\{m�4����َ+П�¿F*	Q�zS�A�r��3W��\R��/q�<Y0��~��	�T]�me���wE���¥u�a�p��>�ʎNN�����B㓵�ᏈC�kS�=�S�>r�V�q���ߊ��Õ(�N�Vzg��=�!���=��?���YÖI �N�*���it�SV�J0��'��+	�dV�.Rq�DlZ/ڹ��Q�=f���1�
Ŝ�z�x��c��#aI�a����"�$?�ᅰ@��foH�q��@3���S�f9l��?��'L(#�dh�������2�6�[}b���c��+����G,^�$�o-�u�������<J~D��YU6��ܙ�|�m�z�	s2��1 �֭@K'�P.�� ��v͞�8�0g#aE��T�ހp���~.�@�$J�Ld���`���j;PA諃
%`�i_>��fob��A���-d�~p��s�"�֪��qb0P����B�^�Fg��7�Րf,��N��̅�?Bk�v&���F�-(c�ג���ti >�
%��m���pr��&�$aY��Ԉ��ݜ�.o.�)��H)dOz'�K_G���Dr��ꇑ?zA����X|P;  �����>r+��Z7W��?���0�KX�54jR������Z��xJy(���NX��i��10��*RPi�ZS���yI���������Y��a5�4C~�Ю���9/�fbO��P�:�so��!�Z�gd~C@%�5�x��|���סK���Ƥ!�b��b����aw��!܇�MZ�N�-������mw�&�/O�׉� ���)�->d����F�KQ:��{ꌟE����ɶa~��ṏ/����¬�3:�W�Q��fU�#�w����9V�/��$�Z�瘎{_ʻ8�<̱Ѹ��YՈ�(�:r�,�t�I��Q�m,�2�4�Y���"�u�)���mLUE�-6u��`����b�g��V@j!�:�t��3b�QG�A�A�aS�O�(ʩ=�w�"����<�=�Ċy��\��v�B�&��g�K�fI̗Rt4�Y�ʖ9a&�Ii k$��JZ�. �D�n!:/��NN�9ȿB�j+g�g=�4V�غ\��Gۦ$��#����DS鰠��/Su<y/�B�W=/����c�_�ͪ���
�O� ��vJ<���)�������*(Ȩ�x�$�|F�İ�q��*i$	����JH"(�>;!�K�}@�*�E{�����N�����e�)�~z��;׮ͣ/r���D�H���J��W=�I�g���,�.��d�>�4�1� dY.�g����l!��di��'� |(��I����Y�|��&��c^g�a̘�W�2lX��h1�[Ֆ��������y�����7DӦ[�cR_�%P���Rai�	Hd���?��i��Ĵκ$QW{_3�p|��co�e��_�x�ۉ!��Uw��b����@���3&R��Po�&Ŕǆ"~ݢ�D;(����k��W�E�9~�	�e6�m�؋���{J��%^���U�iUG,����/�	��/~�i�}�����Q�6J4��m�)߷Pz_��ӷB��~+�����N�|�*��1�,o�_�+��j�����,ߒ�~���Ԏ���UU�?4�9H?����p�d��#E#v�������^r.J�=a-�2m�, 
���A�7l�}?D�@TgC��E�ۺ��-3lnN����y�Ul&#�)%���K��Q��3��-�k���d4p9_U4&k�܁?��s��H���P]���6���s�����S�Sӹ``�R����mD�w恽VL�:<��l�z��	�nWg5����d��^3ɤ�9\��ּ~",�􀘹<?�s�qo�Ej�.[������R4�VF=�g��L��b7͎	�P� n}�ոv��5�iQ��z���쟡�>e���G_�l�<��`����J��9M�鱕'�`��d4~��qaDxE,.�)�4@i�=MR+�I��e��'0���������-K	��� QGN�E�ԥOC���2�����N���6ö�����%�}�5����6�0س��os�Me3�d�!���f嬤��Dp=�GE�d5�����hO���`
�F���7��)Q�g+.{��"�7��L�F�Vn޺]��Z����� Fk�
č��AG=�+s_�'�yS�G�>�@n� �J,��	�@C@��U��'(�l�h;hm�@��h^(��C�YA���h���*�S#Z0��� �|�0�i؀����4kF��?:O������*�v�PsX|.�~��C�4�r#��a���U��|+E�����:c_b,9F�q�wBY���0L��,���9��y���p9q�2�o�\�<�����y�%O5i5�C"�*�U
-l�=�l��X�0@�݁��r#�п�L<�^�˂���<�0�\a�4�iB~�q$$��r�(�JX�W(PT;�́�rV!S���pf�>��M�1��KU�����eT���1
6c^' y��KD��p|�]1m��HɁ��yF'�HF��p�a��S��Ӊ8T,n�a-�u�u춑$���2�wgn�g��G���[��J�J<*��o?�V[6=��Bv��yhtM�/���M�k�:n��R�z&,����s���$8�k̞��B�i�}N�z�c��hx+�͌��G�Zj��H.�6?��Iڻ�d��=!��K8��Ņ`�qO�_2*�x�
�}��hq8�?�]��Q����+�8������3�hC)6�w�[h��,��cj�M���y
ވ�39ɜ���1PTL��DqvҧRXꞖ�0Z�j���m���P\����庤��1���c�hn�v��_��b���ώ�
�>?x��eN!�'��MFY�p!ՉO��3��`��i2��F��Mi�Og����0yL\q��I�B�=��T��\6ԆH���}%����!��2\Gkf�͒3ߔ��\�cT�]S}L�����Id7]�j������c�	�V�\���-�p�stS,ty1�Dk���2�^w����!�DF�
�[R���
j��$3�É�R�,S�5�z�B����)D��例G�L���T�R�|g5{��Ƈ�c �O5�7��>>�ٮ{��)�`n�j�!(Pd�"����1�-��?>XX:��{�o�s�9����A�LR�I��t{XB���y�����8�gN$�`&'wa"|Y�9�m�'z�gw��?�/m�O���i%����V����/�����e3�kٟ) ��a�z0�_��Z����qq�I��f��+�*��S��T��3D+�"��,��c��ȟ��K��m->��F��rpX�r��㺭��e��;e]>���sv������'m�H�����0�]'�i�Z�<���{W�G#�.V3�Z:��Sҙ�Vzsݽ:�J-�v�5եKX������o�cX�jh	�Y11���\<�\����R�1X2]N9w�+ݼ#_Gi�= ��;n�ǰ3ǋ�ށ�B Y6�,]/4q���ͬj#�@5����T�L�:*��4Z'��Ы�'��o��[���su�0���������C��i��e� �L��.q�E�:�����buwH$䅬�?ߜ����P�n���_ч��{�":�`�ӡ6,b�<XU��R������H��3��~� ~��_�xD*�6�*�\t�|�=������gT� 6$C��Xe$b�N�
@)\�f�SF��nхF`|TKPuD@PwL̢��W�RJĀ��v��}������!�t���g��>ǎ.�f��L�M#Ֆ�ː&7L0�nQ~�22�;��
�:P�j��۝Lc�c9�i��yO�<�I��;���S[+���������s\ڀXC�������ָPW���zm���-R�Ŧ,�,��7�X�;@Z�2ϓen�����B�n/\ �M4�C
�V�+���s����ե�3W�|$�
̿��������ڡ\��дY�E��J�5O���"��\\V��R��9��@����-֓��̈J-��ru��OcNoD�[��-��Yʂ��,��B̙p�����i�`*9��gM�J1�1WҔ9�t����m����%�^���P�7�R�w*@ږ�ý'!�'�t��!z����PB"�Y�Fb�)g�AW����<����5rx�y��P�RX5�g���u=q/�ܠ���W_VR'h��r�\yYoɧP�Ko���U��\3���gR���&~
+|F�K�fD���W�
`�N2�x����H�w'$£��Gl!x�)?�(R5� ����)��
�9M�Hy�N�O�e��[`apC�|�r$�P�%���n�oB �u�Z��*I�:��bќ!��n6���.�)	�`���RQ!ª���N��D�ay�7�#�;]칠1���.Ϊ�M`�mV�FQ`'���V+Ce+���Q����@U����e U��&��Ly2����[f
�H��=�kYk)���bm�63();�� ?��AS�,a&��&�� +j�uq��XNq_Q$��wQ������'P[�j>�����c�zb���$gd��miVnɡ�G���B�&ގ��<K��gFټD����^���k�=��C�.��׃�c)"�	d)"I$UH/�`Wo}jL=�g�����)�aW�r�����Hc�V�y���?4M�^l^49��{Ogy\حm�: �+���L��B:���h9������PSP1\i�庞�6j��i��8{���
����y�1��Z�[��4���3;�h��ȹl B͌)�2�6]�S�F��v�?�k���*��Ƥ�N<!��<���63�+����g��J\D�}�/1���Q�/(Y�T�)�J+��I������\���B.i<얝%�� @t�ն�~ե�2L�E��!�?��	�B��Vq

w��cs����4�寘�)��q��>�Oݐq11���6V&w�Y��9�O�+��M��N�9���hH�?z���P�wEj8��Ѥ�T��E��K�h�h><��!�!ZW, ��.7��DOw���9���_������g<#�z�ї����p�,�pE]�A'�Ky����D����$�]�|�Qʏ��~�z:�G�5�2�#L���G5TF�@�����c~�!���6ِڞx�w]s�D�w�c$�%�OD��NcI��	�(���4L)�&�z��D�̪�=��[�J�N�����'&~p�x��qn/�� ���Dq��4-�������|�b��[BP:m?Yq�Xm��8�r c�.��V��]�F:EfA��>BU~wq��9� X��ZJ�{k��s�e%v�Y��z"=�����ޚFBj��{dj��@��չ]�q��R�b�E5y���J�aT9���sg�@�pړ�S��DĴ��	���GȬ�N�3Tf����F�qA�-��l�?i���f��i�5���mT�L~�G��A�7�>��C�]����	�ؚ�zVN�1c���x����������3� �Sb/Ŗ;f�e�xRnr��"�ؑ`���z8��w:�͛n�M�h=P�\�$��a!E���C(�Ef���z���KO���
H�)�oe��\��L���+¡N�"��#'r��Ō��!H~�������$�̄�,�� ����w��� +u8d��T�e=`㥩=\|%Eh��M	��.D�H5�Ʈ^���X����\ ��ž�ؿ��X>)�\(,�sU��oV��3���)ͺ�٦H�'F����.ፄ���F���(ۖ��� $Ɏ�x��B|���8JH�J�������W�H����`��)��'���F�.���|����}��n��?���|�����ezY�ر��٤���>q츐j���0*Ǿ�������xG�i���3"�U���j�γo^ �޶y�^c@��+TB��v��a�@c��Y'���psו��8���p��<E%��bm��P�F�*�$�=	�����ˣ �.���0Q�[V��e�'�����H�kq�E��H2�������{]I�1KQ���?K�+9��G˪�-���fU.�D�c��i�+�o���U��P����h��4��; �5Z`��v��:�e%-�'wQ��א�fס���͝�� r�R6�������	�,�> [´�Tw�(�?�
�lP�*���gG-7[n��w�(�������G#�s��t�@ޙEB�J���F��1�$�/ǂ�<��ӗ+jՈN���-�nS�%���sj�jE��+V���77vI�A�~����D�ޑ�;�<��ͩ쿤�_�W�/�&uG�&���i[iA78��B5����Z/o�*���D�V�����/7s4�nr'�W�RTj�u���i�#��ū�U�*6!� M����iO	<O!N&5��e� +�#����A�?�Ы.P
��gęf��]����̷L�#��[	��,�������.������+�8�\zNO����$??hǤc���k-�:͗�=?�wԌ���[3.���!���������St�:Av��Ӧ�.v*B�/}��<T��	�����V���M �������F���3�Fp�J��4D����L�I4^!�ԝ䳊v�ԌE���c!��/|G����
v�d%S�DH��ˤ �*�za�!��a�}S1��/��#��v��G%�f��=�0��o�*n��r���d�cy�0za
X@�xn
l'�)�2ڎ���T�d�h��6$J:B6װ͏M��Ad1�;��}U�M���-w"
�pef�%�������#R���z�4�QdG��.� �2H����}�8���|��U6��`�!�����rr��U���=��J;��_�AHh��7���gcuG1�C��
��4�m�����e$O��'X�{X�^���^���_l�"��K�>u݉q��>�x���k���ç��eZ��t�g�{�
 $���С����.}c�Rb"m_�+ꡖxh�Cv&���,�R�\�����^{�hb�Y��D	/w.�g�8K��MB���顉r������]��A����W�ԗ�L�n�#�(�r=I�誢���%���1�~0�~���~Ƿ2�hѳ�U�`X���4�3����8Ge�XN�0]�.e(�V�WT�ob����j�M���wGx��R��8��wX;�����=z��
�Le�X�]0��)�<���0EL�2If�M�����]A4L4t�a��=�<��ؽ�R��Gbm�M���I�5)��=jg4��G�֒����6���I���|�#řZ]9U� ����Y��ܾ�ƒ���=R�<���3����(�� <Y.�)�~B����$���t�	鴸��.l�'�l�����6,���z�������6t�BlJqt��?tF\�1��n!44�Ӷ1���g�c�����/�<������e.�F~^��6�N����h�Y�D��id䌏�.YoA-���IL�$� R>�B��#8���<����T�ۂ�M��{�Ŭ�PQ��%l�%PԀ@��AƁ�ZٲYQ#�7[�����:|�]���H�u�.2`�Hc@�H�Q�F��Gr�����ޔ�^҉��T��@Q�i��`�{�d�3��.��l���vN�xV���&s���6��S��ax��+(�?v�DJlV�:��%hM�yo~�T'g�jj�3L�|Af���,w��"]=ˇ��AMkI�@�@�PV:���_/=�3JK�h�)��%uş�M�ǶͤN�����|0�;{���0`�9�����v���91=��i�%�j �w��DB�M�xP�e��P�V��N͒,\Ǡ��ܵ��KXԘs��d��E����6|�c�s��&O�X! �`r.�`V��<���`��~��]c�)hJQd�Z !d�Y5�;3��zո�+�-^�|��!���֣������Î�K����O����g�����Gx~,��΄v�^"��4;k��n6�O�T��>3�xs�KE�$�{�[RP�#N�L'ݿ۷�i�8t����1f1��}����lM=*;�a:\ձ\�5U���->k�kӠ�q��aue��'M��/��ԓ���i1U)����+�Pb� ���Ac����o�W�L����³��RV"H9�WN}���&�	��ͫ��s;�|��;�c��p���:�!w�]y�ql�����C�c��ti?`�V_�I�'�6h�u����۠��WN�ʶm7DB(�/8���Գ�f,����\�t.Y\���m����<)�^�]w�����@C�r��;��֛e�2빲
S���w��^l�ed;s�3҅� �4�Ui,�����r�9μ���\�#x4��ٷ����s]�G���H�9^�f\(��g��`܎�r����>�4��7�tѪ��ܕ�ę:��sykh��a�T�����*�����
�Q=ú�x��dT����1�&#�0�nz��q��B,}�/+d	��Eq�����y�t%0�O�����ְ"���oJd׻Z���c�.D�=����RIG��-�Fmf��p)8�DU-�=ܣ��9�u~˳)����ǂ�����9�G���G0�<D�wLJ`�����N��K�]XN�׶g�D�Os��_a���į��eČB�;L�a����lFO" �B��f���AC��7�	w{{+��?l����y��:
�>��Ӯ�����/�$��:��5��,w|���5��,���*ђ���I,k6�8���aO�F�xh��g���L��5�>�s��f�����h����ܺ���$kS6�u�����cK�m�1�S�5�D#��j�W�����?7,���*�P�X�����J�&�����7�Lqeo{���s�8�a�&=�}g���%F\��M�)�E�sF}�@�c#_���v��ܵ��P�8Z��	V2�ȟ��i�2��� B��3�7�d)z�(:�[��������n�n�䧽N~Z$&A�_B>=r���~p߬��k�_�̕ `��w��p=w�ԏ��+�J�<�֡�z�v@Ǩ�h5�^�I���G�P�(��5��E��4>��pX��� O��Ţ�	��d��Π��>z�����������	S��h�MQ�땥��ҡX�3�-F�s�����~aC�Xt��������6
nFxy^*�a��/�R�b<��»\�@2ͣldw����ۘD�N��;a��K}���~�@���8�~>"My���(X�{�͢�M/#ݓV�M�ء����j���ff�.�{�����s� �R@q�c�g]�"���flp��ͪ�f�>���U^�0������L�u,X��8�/oi������.�`����DƧ&���02v+�t&����@���={��ʗ�o/P�'�`�&;��G��J�<�O���O> �δ:��7��n��f��k��A����5�kf׸�-�����'�cL̒}�������P�3e�{qx����y%u �������S�)��cM�O����݌�Vk���q�_+vt囇���y����K�Fm���%3����`F�l�`�K��j`Y����G�[�"��R�aF(��|4<��\�~�apa�$W�ݘD�����0Y�Hko=�Mdתּ�&�O�j`�x�.@����o_�����d�4�a�������"��Xl(�����z�^�I�?LV�f/d��`�9���=�F�{�\ʿ}���~���{���x'�I��wP��)�k�û���� (¸�[�X6�=��1�.�;4�U�b�����Vdg����$?dOcK�0�b�k%�+�D�ALo�J18�I1+�+4s'� N�i��Ju y�/�%�(r�ǟ�s����B
�+�$��Қ:���?M�T�cy���uttaD�=ԋ�y���w
��b��w��jp����Y^`?��+�X��f2��+����V���,e�wx�S�ӽN\֜D���h�3D�v�M�՛|2?Kil'���Ur������p��Լ%2zj_�Gk�f7�9���b{Ɇ��ڮ3k�W��l�#p���xfz;̏��rD^����<!W��[I���b�L~(��3�GCC��;Pd��侮O��s��[<J���F��
�i��6S����ڵ!�|�E�dc'���  9D"H:���\�i�YOUI<��D
S�At"�̡�VW�EOU���l>"� �����3��K�a�9APΙ��e�:�L��0A7rx��V�U���@Q�sʔ�����B�hrHS��i���.�Kܴ 䖧+4�-�L�2��!��
�܌�d��E�	�ly��9ߠ9&5ewŹ��bb��������3 ��  �i���r�����>����X��8��:Y@�XNZ���iO�Qz���Z+�g:�V���Y����RO�TO�;a
y�M{}}�N0<��F��l3Ωo*�\M�v[�'#2ˬ989 �=N�pa9K�Z��_���Ofb�����3����3�U��>�������}��&����x�d������-m�]i�v6>1�@s+���)<�ar��^=Z��h`l�L&g{�qv�[$�VzV���th&2i���4���_C���P�c�.�Kk�{�&��Q �Dk�Wo���[p
�>�Cn��xs��)Q,��ށ���l�*��л�߼)�Ζt`@��#��O��Q��wE��APT�_@y֮��P+~�~��|Ӟ&1���0I�c��R#̞ ����Cyd��)�;�F)��c#��n�c>���z�v�/; �h����և�W�s���y�U]-���NL����HE#y3��<�zpIG���Bxa��,���D�g
��]�usu���p���a~zzj�-1 ?S�EhP����YRO��^���^0����쎎$��"����y������x�0�V��S��a���m���U�-��]��L������OY(oV�Y����8�c�X�i�i��Pٱ�� ���*HX��̓@�C,�<��۰�	�t����a��>+��f�e~hr�M��Q�:s�ƥ<O�-.E+4΢P����m����A��L��^�p�c��l��hOH���À������رa��O��c�ѪwA������?��apX����[���QT�����h�d~5u˗s]7�Gf��w��<���4�0�A�D&�a|y�s�:��&Ɓ��ԋ�f��P!'M5'�5Fg	��GD�v��.δ�]��{y�+���K��M&����E�F>��E2���tO�'����~	�Av��F��'S�l*xz���͠�ݱN�	B�k�B���7�"Z% �4�K~�v��x�-���X@��s �T�8��Ł䩬:�j��C.��@��k�'�V�a���<?'PS
܏y̱�3���
�
�
�~���'�kQa��@�)�ᅞ3��Q�zeg�x�����P��h�E jk-Zʖ��f��I�W��/�=��м��y*�����C�g����l�[^�����ZO<�ʦ+T���נ��9'�o��XR��y<!�YX���7 �3�	}"�<a(�K����]Cl>��xo�}�
²3ړ�G�S:���o���6�s�@�׋4B5�l6Ȼ����yت[��(�RT��ü��{skZ��4�L�P	�ײ+������zm���Вn0�	���W��8��GK�vf��Q�Z&S��=���%�����Qϛ�I�[Pܩ�aO�̕)ڰWv�oh�%�&��C��fY�:}���_R��6tqt1�}�������D������R*g��yJԵr\�75��a'���O4>6s_�]Z��d�p���S܆�f�J��" ''�Q�ڨ��b�Яr�o�,�79u.q��c[��$ͺϋCk�����@q57}V�ۚ&Z ;6��48�x�LT�/�D`�2W"1TO�KS)�'ʅ��K!'~B��S��{��G��AM����#�N[/qH�Ϥw����%��#���� A���b'���km2��<m��ʜ�j��
6A ���QWU�����3�n���aR�	Z�D,z�q�#ٖ<In���A�ݯ�M�B^T�qCCh���g�����S�<�z��c~jz������
#2�����"Y�(������2�fZ[�|��؇i0�X(�'t���\.l��iP�'}\?��TZ��D"Sd��	�8;i[F��D凙���X�,�zн�U�����ٝbT��Sit��5�^(z��A6B����� T� A|g�������۔T�7"}�A����q�~Qg�K�VZ{��^��r$���r�3��U�tu;�/�8ʴ�kBn��*ʚO�C����`]�_�y�4cl4,�hR������;�ZGpBJ�ʳs{1G��%>d$���+�	K����}�AɅo<
v\HԱ�^K7���M���ݧa�e$�� >l%�)�+�b�u�4�v}8:��:
���0�9�mH���3b�&�g��]N���������D��F=�5h��'��(!�L��k̞�*wP%��϶H`Gd%�������)���2�iή?PJwj���f!�y�%�
�
8��� Ƒ���Z��/_0Z;������԰\������h[��s���J�h^�o��.��_��=D�bN�Ȭ6�=�Av�%�i��m�G�(�e�5�/�.�hF��16�U�:#��)#سco�W{�E	���^�1R`O���`n�\�G!����ۈX������( m���{^��̴�ut��!o��+Uߺ��S����@@�L
�V�'nTI��J��~-q0�~��	�!~��J-h/�Nۋ>D̤��h'G��j���M�OA�t�������7�ХQ�
��2*����q��b�R0�6��O��Oy ��Tq����(���7g�T��h��Al�G��*~�02���$�=��� �)�<���D��jWS���cy</'�d�=�]e�|\��r$�@Qu60�q2Li���:p��o�~ܥR>�4>@�&ZO��S3O�u�K3�zN������Թ��QN��/�I61�K hW�>H"�%�:���	>m_U���뵽��:��w-�#��غp��F�I�^wF@)N�u�E4<#Q�2T/�FӏT�}�ě�#��{��[����YAKi-���h��=�@�[��ki,>�dŭ�>��N�I\���0��u� %��m��F�o�w�LG�<?2guYҰv�˺ӶD�0�}z�'�M�ލ�+�b2����3s˒yV�B3q*��E�$������c��t q����2��2C����.�s�A�`?yB���"��児�H��"#%�`f�ca܉�e��r<K0Zi����t��*M�1�����[��"�=��Z��z�����7���-����O�g�0�k�'����ĮΚ�t
<��QSbׅ	�c����4MZ%MZ�3G`�@�%��k헱�8g�� y���^�^@���@MT�n{.U�m�Ety|��s����r�żN���!v�a��i1n�s�h�����r��9I�(���1߯t��c)p�*lAճ���������{�M]1�,�N+�TD�?�<�]lƆCk�q�^i,��j���t�q�؆��b�5U8ߌ����-�<RW��'�D���P���=F��l�'$�ꣁ��5peQ�i�,���n�A����*�����^���ZȪ;5�lu�T��ӧ/�כ/��t �ZQs���%R��b�n�/��w��a���n��w�puy�}<1�rs����3�|�v'B�{g��V�b3�3Ա͚�*��5v�`=��ůwiq��F/�[&�LsZ��h�;�֕�w���E� ĬGb����k�������߿c�3�ڡ��\�&�_h��D�ڤ��A�A�a��Qخ�Ҡ�F��p���Ԓ�{;���# ��ӣߏW�m"�>Bʞ3��U�
�Ѥ������`F޸�ǉ�h+\�`ĞS��?ԠP~��X�H$ӡ����ƻ�3s
^���D��crè��&����c�ɣ,���� ,�2��E�G��{M����zYZ�㵝���h��M�2B��$���u�B�=�A#~��ŧP'������7Gbf���Ѧ2�������n/��4�=����s��5�%PJuE�	��r�@Wh6~k�o�_����?�����P�t�����HȲY�Š��Ь&�(fù�q���,�f_&�%�S>	�a���G'���UBd3�A�3V��߯�
��>�-����c}(���7|s�r.���1�c��rHUP��������_����/E��qR ��	��JNxn!Sy'�o2��X�b|���ſ�H*���0kwB�L<{���C���?Hw�AI�A�%��� �ōx;�6�n�]M}�5�V���aa�B.k���7�0rN���9#�p#��\_�OX_s�\u�2c%!�I09 ��˫���x��$�PP�A��8A�{J���ɓ�"|n������-P?�}�h�'�^�7p�#R�;k/$N_��*Pf��R���/����G48� ��{4; s]@Fd!��."��m|͡k�)����>jdi+!x��Ъ��<��P��,��Z&�@��G��R�=�� {p.P�׈}�������]�)�g{�����^o���C:�ݰ��̮����kU�����?�$$�LO��+.
��d՜D�t=g��
@� �8�@�_ը��Q΂2$�f3��vHs�t�Eg��9�+����p���Tfvp}�ZS�ᓅ6ZT��g�AN�Q�ة�?L��-�+eQD�<ڢ���!��c��B�܂7K��{��<5>��Å�^1Rt�Mr'��%��H����v^����`�^�����L쵷/	I��GPު�ő����J%�i���)$L��U(Pzzoa�491[�@�9I��ޛ���a�g�8w�3w�
x'b.�Eh��D����N�s�u�p!��-a.���r�������Iy¬_o�e]�-���Q�;H��)��)3ʎ��{L��M��+���o���g�h{&�^{�; &��*T�M�Ü��ڌ�n�i��S%���ΐ�0w<��Gz��:�S2B#LԿ�w���p�����Q��gM`7b[�ū� ��	�=��t�CNҷPJ��o&����Ȃ��F7��+�7�C@e�6�u��A3���y��3�jH�&���K��y������v�*|���˽�)Z^�(:�hU�����u` F�a��+O]�g	;��b�N>[5�e��	�Tj�@��lG��Dv���*~��ߠ�sf��ȉ�k���m����\�y"�ϛ��S����N�N����g�?�V���4�c��,���.�mؕ����Φ8�#J)P��Sg�`>�8�u�N�QzN��4{1��+w��4�-P�����x�"^w傰{�'�Dm<53@F@�"�Ѯ~|��i*��Gk���tDpNgSxv�,/y�%nOW�ci��t������%�����c�x���y��f?T�V�06�Q�w�q����e=� ����E�_��&t	Gh�%c���+z\FM/��³��:G����$��P���j���0��F{�W];�7��N���{����*n��<�ızѓC�$�/N����|����Htګ`I�թ�a��T^���8��\]֎Mr�{����i�R�m��9�G��_����Ix���Y��j��h�*�
�T�ݕ�|�Cv�ւ���j���1�B��fpN�*նS
��k�r�T� �DOʋ'U�`�]/�%5j�c������3�?���Co�9�q�I�/7��ǫȇy1{�g��)'9nL`M�E]��	oK�7(����/N������5���_��J�Om������u�� ��$�Fg���0V��=�����5���bc�����w�R~��8v���1֍�	3��WC��-�n�$�ȄEvL 6�������(����:��zYW:|�j*� ��ڼ����orOm�6��\�&���\06yБN�
pn*ȣP�ނ��׼&o[2�GD0��ؕ��Rݱ��%JĘ�\xi���ߩ�b���?}�9�)a��* ��i�lgd����ACP�Dc-cAi:-#�:,�h�� Q�;��9�e���tR���+c���nf��\�KC
Qک�9������׌jU]�<dcp$���� �����!�$b6	��隧.N�4�[sݫ�`%�{b���*����=ξ(�b�dr�1��CV�1&4�`�b�F*<��>˛��9�I�_�_���n���̬�>��Я^��55G�B�̟��U���v6����������B��b9�
�`���j8/ D�����RL�lEa��fk��Hݖ/��Ym�/SFX�W,�6���&)�G�fl��RT������]T������7d�y���jf���S�vr���p#�g�#}��UoA�pb��o8�*q �/l�y;��F�7?���Gn����_�=�)P'taqf�d�Y�,�w?�����Y�Fň@JR8��.vu�?\;z.�^wK�A�0���\��A��F��J��X�#?�R�;��b`ѳ��? QP�����B0�/�2�}�43�����6���Z����ҿz<� �kA��7ҍZ;D��*`ؼ��Z��37�H�P��5sk;��YW�j 0t�jI���tr'�Is)D`b&�~ܮd�_�cx�T��	Y��x-R����4�'���� )�n�oi,%[�����99?��[N���	&����5S�o۝ō���!nA�4w@������POx�"U>�c�E|���ox�)7�W������hE��;�ԙ��y[�U��,v�v�gSG�"����?Cq�JǱDz��U���œ�8m�,�0)?Z��^P�w�>?^r��2B`��̭��bn�q� �v|7���.Tm�*C4�7��A�˽�:M B#[,GU!!205�7]F����/��&�����[	�+5�#2A�p�c��5x����?���|���gjs܃��df�7M<�f �O����t��);�yI�$�"	�$�jƙd��:Â����$T�xGs��d��ߋ9U��܃�3�*�=�����4N,�s�� ��@�bM���ɸ��(��ƙ04�Z�f:Y_�2�������5m��5�x6L#RP���0��1�Ӽ���s�F���6��*w��ZtpصS_KMdx�D��[���>[	SDp�u���4ɢc]�Z������v=��%.�7-DZ���S�_]����ݚ]t�K���C#��;f6X ��CR�{��Z��7��-�`s?S:�� o�~�S�%0Z%C#5�vD�� �I��?�T���J�w�|��7��8�<z�#��d�?/i�׻^P��m��=��{���>�A�I�xw�1��p۞���x��k��L)��V��,���R���S�?<�h �UӘ�h�*�S�$48 ����v���f������#�К�1�Z "_�Zk.Ϧ�da0s���h5�@,pyy���ɦR��=�s����Z�h��Ą%�*,��w
�B��a�J	IT���������+�Q���M��CSn�hI��q [&$x������h�> ��%<�ƋH�N��ǬpnC#5<'�����W��JlF�n�[5���`�� #�p��_��߭o;4�G���4�~x�$�ެ�
�Jm ˟� �����Ţ:�Ĺ6��Ȼ��m���� �\�k���l�L"��lz��-?
N���$�?�����.>��TFOV�Hsg=��ᜄ�p�ZS�X9&��Ύ��6���)L���:@H�I�������d�tm�]��S�"a���CP1=���+�ލV\�b���7����2ۦEZ�_�����G��Ӧ�Z��=�-^�餕u��)�,�I��uss�xT�Ì=��O�H�L�ڭb=��u���gX^a�a��i�WE净;�z��[�m_g�0�_��0w8�)+���+�>�v�71��Nϯ �f�b�\��ґ����������B��-wVz�5��!Z2Ҩ����H((���P��ʬ��cc,����kG��#U�)�]�W}��"���.��$��;q�|�Mwɓz��~;�H���0�R��a��v
�&��^�V����C��)��$g�R�$��)�E�tE�`	OB�A�i���x!�ܖ:0/G��Y��9��߅۽�s.=�qK�"Q��u�)�aiXG�����B������|N`���� [Ԏ�ǁ6H�P��7%�$���P��[����HFQM0C�vqC`Hn�aѨ�����i�^P	�U�@��T�ö{!�@W1�(�*Uy+���bb��HuE7-w54X�d��WGvae�n�L��c^�z���-�~G�"|2�+�qρEĢ�`���h�ڊ`L�s��^��I�=��g;@#�HUN���(�+�i���(�uG��;�MQ7넶�w�'�ĘV��!���\�{s�]�Hc��H�p�D�$ɿ����f������W$�%������fG�ٟ�7�;�<NP\k�dZ����y���}�T#h��o09{r�����By�5��j�SB1PO7�?��~�8��be��T55iŽ�A�� �6���ՠ��ұ9�i/�D�%�l�S�ҙ�)��@�x�l��Ej�s&����P�'���7Eml�1\����X1�}��v"����b�(d3�K�y�t����6hJ��{�1��ś�]"�a��������,qB��K��;���e�(@���@/l�Z�@
H'xT���.PsQ�H����rI�F�`f�ǒ%�q�uT4bD�i��)hf.����
@����J$�/|_ߴA�Z��_�1�O� P7���M�z�Τ�h��X&;��ةH������TG;�wfő�>$�
�rI0W"1p��K�A`�:��^��%�ut=��/y�i��9L�o���"~���`C��f�])@1dUr��W�L=��\c�˲���C_�V����l�}�@i�4�-�F�Z�(�x��'\����\��O�/ϑ��켛�kg0u�U�uO�+)�pf��h�Z��R"&�J=q�!.I���n�ؕg��ˢ�6�����r��s����s�%�����8עSwDq�J����S��o�b�ʆ���4�c�8$���m�3 nQ�X�!����J���iG��Rr_�F�Eۚ�MB�p��4%�p"���8���yh@S:W�"Ɋ=��	�#�I3%��UV7{��NTgR���;��O��j(��v/uJ�tFn�`'�o��Oº+2��ʛ�w�no��MCH�Z�)���&9Ӥ��W�A$ܽ�痯ym2�4K#��p-��.:��%��n1��J�'ކ�C����:5��%�>�(���o����tij����6���u�	��*3�9��'�ײ)�lV2���&�4�B�8r��,N���E�uj�җyʧ��-n�ȯ�r��r�6��l������fr����4��%zv.��6����c�����٧�o�4��c�a,)n����|�
�ڣs�����	 4^�G�?�{���IB^��L���mݒ�������wWJ��4�ȯ��R��o�Ǟ}��)�ߓ>��6P�?���K�#��"[^|�bOM� �8�7�A�<y�X &�(V*]^�!$���3�g�+5�;��F�b�lT�&Ǻe��b@㷯�8Q˚��ڀ���� ��ɪ'Ӥ��2��M���v��q��J�
�ϥR_�J���*���,;ǃ?�J�t�G��4�w�O�.�0�x�[ c�y��<��ȍ��)�'��t��3 �oXK}�ڑ�O�9w����t/У9~��^��ػN�s&\:5�cn�pZ�=��ݒ�O�y��F�5h�,��r�.%�)�E=�|�TN�u����O1�B0Ku���RS����_(g]�1�k��[�_��V�^��7���w?.�@Q�������,Q(�9�B�Jw�/̻+��u���2�55hfv�G��_�k��m.���"�!�C�4�_+گ<��p�N{�x(�B	h�֤��%��Åfu�v��8^�a]�N-�-�*%&\Z��1��LQzi��X��QI��,(`b�d�B.�so:Zq��p��riM�g^^�����bg���_q9�n~����(�#�\Fz�.g�X��
�C+b�z�wU�$(,"K��6�e6�SVT��sӍ#�-�~��L�WV�J�ZY�V�o\%���1!�e�ZUʕ5��4^ҥ�
