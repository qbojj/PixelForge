��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����P�^�Mqap)%t�?�&�Z�K�*���~O��in�ÇZ2���RG����R����k:�H���QNOR| ^{Ua��M��m�:�$���/�s�~J{]������oٽ�/)��R,�9�Սع�T��̈́�ͧ���NW����[�R����i�IB�z���6����e����yv��\��e!���_Z����j��E�i*�!�&�v��X�'��EJJ��
�u��|A��O.���ۀ�S*����{2�U�R�i��];E&|��$�d�ހ���LJ�<�[�'��r�I�N�֧=�H*�(����դ0�0,D�Xht��s�3G���[b-4�i/Ke�cU��`��ă���M���~R��j_a?y	A��h��fpLw����#͟��,=׬~�D�js�5|��,u8�̨q��F�v*;i�*�.�ܭAȑC�h�#�x�F�#�'Ϧ�=��Ι��Z��3H�9,�[�5��4Be�@�+ө}a���f�0!��8�_��.��A�WZ��w؝I�&S/5J0�~J�Ո8GM;��4�8���.�Edk�����W��Ը������f����ޔ[�I��g8G5N"p��To�շ<?��i��z*�_�u�����#	��Ԏlmm�����Ԋ���#E�~'&HG�_��3�����!���n���I�>O	�$E�k>��4\�A���X�C��)��];��,�'���Li�|��vB+��:e���D4E�T@��s��ڿ%T��i*���/I�답n�c�kӃ��KV| ��<�ʦ�.������4ˠ�-Ys�'O�����~���>���!�b�^���q��ZJX�HՄ�i�MQ��F��7o���r��i���� �ֽ-�o���K�@��ľ'_	�]��m��Gv���:Q��T;��NMl�_���z�f�����7s��Ѡ��upX�,���$� B9�O9L�q���Z^� �)�<�����"y���t=�h�|,=��U	��KY�k]k�;r��]��ͩ>Db���+\/(�SS���a�)'&��������vc� �*����S�r���q�������	?��շZmB�Y�e�O�Y`�-*�Z��8jz����G45�cx��(�̯ ,�4��D��\��*�Ġ!6�������.�۟I�P��$�G5N�H���c<0�4|Dmq$���=�����]�Z��qݲ�4:P�X�}�"�����t$Fv�R��H��GзӜ$��I����N�p��^�������g��5W��)������,0�3��� `m�[|Ћ��H3c��R!��}���/�2CK��@�j�p���
��׫L�;8�lElCQ5�fn�#]�MXW.�S���u��oD���R$G���	���OH�		}+�������w؝%�ф��{545��C�Mڻ�<�*xP��hO��Za�M>kP���v`��pw�Jp�[Ȅ��k��+��6�c�m�E�w[����
�X!��3;{:$v�G��m������7z��L�R����ؕ�W*G�p�v�-|���yuЊX��K����C?��%�l��3���I�׽f����^ĬRu4�M<[Z��[����P��s1Z�݁����-�W󙀊��>�g� ;K^��U�!e���w $�����d�ލ� �Tf#@���cӚ��.��y���6kw���� ѿ�89b�l�8�����]I̎��T\���fƑ]s��u��8�)�k�=���gC0ʁA��a�Ov!���@X�x	\Oz�J
Ls��:�0ֿ��qaB���Qa�|�6S��|���_���:=ɔ��O�O�b����R�b}e�..ݥ����|g?'Gg�Zm\��C����Z����*��r�ݧjP��T=���6gM��y��1V��dnډ�:���%�S[�ro����4���z&V��)��K��Ff�B%u�����>�D��hЋ�.ur�Wk�.�p|q�:�?�˞I�s&������:�:3UZ��xy�qtƿ�����R&���u������Vu�(d�M�-*����^"���A��9J=>e�����5Q1)��qۏ��r*�ы�=mui]��U�%�����
�j�OJ�.��W�A!��$㕏U�w�d��4nR�H��'%S�Cr��D4��GT�p�1���NT�d	�7B!p��vq$3�²``�mH�DA���4�?|3Lm�F��k��/�b��L��K
�fP=�e|�����!����Rl�������_� $��P������O�1��gN{��49�
6|+[kY|J5}%��R�녧������f�^��/c2I�7�v��TU��U�%�)���LݪU�;�5�
������'gz��.O��J��uA��9��],ŏ����*��W����.m��8���������	P?$�[�W4q�7۾S�\�dp�������	�F�w2�s��S�!���p�)�;���4��I�����o�z�F�W
<�mY�ڎR��.�l�F��E�A鍁~�}==A!�4��Ę�c93��)����	�Ih;��f���-��d@)1�%�0��ڰk�'���BZ�3���VmU�:�ތ��Cp�c
����A�8Ka�<���uz�ʢ��=H��6�=S5(��(zq�헯*�w�q@V���E`���蚋�I����Yڴ�MP9e�eE�.�����sy���,�r!>�-M)]���L i�����'w���=�����0���Oc���c��b��~C'<��"��<��KNLL�H3�� �BNp�f@*�@�KڔDǀM��#��Bi���X����,����g�pX���%��[l�1���xک����͙�,#+`�^ʼ�A��\_߅�;!(�/o:�be[OL�Bb�GX�:�"�A#h-}�Z:�gMgPR�'	�0�Z��^O�ߏ�Ϳ�&a�W6j�~�#��+{J=�
J�G��X�Q�a����١{H/�+��&M�Ɋ�XuEYjՀ��TXN�شn7����5b��聝nhV?U�O�K�1�+��]*�pX���E6��FS��A
^C/�q'� NS�_��qۗ�!Z�p���������F��FE?0L�1�����	��6uC�E�H;��(�[)R�B��Ɠ�7T���I/��M�)s����%��wJ��
�d�s��h��W@?SӍ��(�l�|���`>��ĮH��Q�=~R�uò��ua8|�W:���2�YN�֔	{E�l$�K�&���"Z��|��<a'�t8��B.뙰f�Y5`�S������.K�,'�72邟��eg�ld�>Yґ �Cn����K��r��w p���Դ��{|·�*��,v�gVߟZ��8�I ��;ݣt{�	��?&������5��- ZH��<�#�^t`Wy��XB�Y �5Eq�1l}ql�ԹH$7&�Fp,l���B�~�q��q0��25;O?��}�녙���`�}u�2
�%��ܸ����'���,U5����|8������Zp�y�T�b�6�vW�OO���P�PH$�����s`��%� dkk��[�g�'Xx��ߦA�����u{_Y�h�]���W�����$�Ƀ;��D�3��-�u
^Dq�9��$�2�gR����M�4mi��B���6n�=1�fr�I˩V�����MN��=�6�'EQg����ϖ��e����I�j�	���/�����*݊3����uwC7`�t�KkfO,4a���>!�C�B7���ӫ� m@��몃�H�u�n!âx"mF�m%�ZF	����i��CJ��w,����q�=� ����+���)�re���QJ��|	�5�rٚ��RW���2��d�.쀮D?Fr5�$?@�Ҿ���ҩ:u-�r���yo?���C��Bu+ٮ���']`�~�d?�J��#o�����&� _0��*6�qܰ'�-���y[�گǸ��P��r��0�bz6Jk�-�]>�9����B���ЭQ%M���m��m����1����-#@~j�3Ѕ�@#_��ڄg�eе9,��'��H{�P�^��x����L:5I����N4;4��s�?��q�z�n(��������}�%���%QImWe!!�H�L��3-Tep���ж�(I(m�^5�q�!�я}yE����]�0s$�/�tm=���w���6)XL�l38}��d���>af"�Қ�jۜ,��p�z���J. �a0j��0.%��9�굧{jP�
F|F��^�q[�׳�Uj��;M�������0��N=x͚���
��
���e�mD~C
xq+(����oP"BCCN�5�t��z��.6{��>��[7�W��ȅ%�
�9)�ja���\RS�ɊK��vZtb���6��ѾOg��|��BHa�rDY�q�<��Q���Ob�y+`��9|U���a�E���
�ʔ-�+��1I~�L�O�:��dw���v(Cw���-2&�"�nQ����ܝ���x-rY�Է�8�?�^���Х�nL^��.~G�uW��8���A;@�{�i��%�c��؎Ms%�$��'���l���K���շv�[h"�q%�\oC7F׏{q��������.�{�ɱ�뷙ٴ�77��5%�<
��uJı&�H�T�i��C��TƦAq�	��ҳ��l����8��d�U��cU*��C�� C�����d�/���cEǚ�rڃi�n��4o����G1Z�����1xU����m�>���|�1��\9�AS�%�8���1������t�=�O�2��Yu��Sz�Z�gCL7i	x+�c�.�	a�����e�,ϻ�D���_+/`~2Y%x.A�c��I���礱gF��	�ik,��3��x?�Z��YVPSm[����������2���/>�ȥg�ۧ�*��WV��d"����Cq�W:f��U���8n'�\1[��O��#�Ŧ��Z��3�~����6V��]&��8Fܸ	��.
t��Էe7�iD)zk�ȟ�H6Д'S����r��i_���{&�$q��5�ak�[?*"l�~�;|s}�8v��@�dLѤ�>ey�<4�+�	r�,�b���^r���^����<�UҡLwY�T�t��t0��`���	�T�B���%AҬ������l�X�pH슼�d���s7N��?6�Q��ވ�{����fP=�'��N�kQ�4��oa\�8D�W�<{���n�_e`k�S̸�ȖB-N��6؂�F�P�����n�/�inT��i�˾��$�$K���ʄ��6E�|�� ��f��yJ,��*M���6a��o0�r����ٴ� 0S� q�s�V��H��h��4� Q���/���g/�����1E�o`b,x�k�k1됐9�X���v&r�Q���J	�0K�['���ʎxv�5b�%Rݏ.�@4��%�v*���N���4�ze�����l���(~�~������}u� �6�p�9^�����nl�>�ak��L���=H��PU��CL�!�u�'�fy|l�G�W	n��;�6B5gٽb�o�%��Q4�G�tw�̬q�jkX;�6t�[�R<�����@1hi�t��3MmA@g�0�"�gI�Y���:2���n�4pФ�v`C�hG�l3<��"�P���|��=��4JZ@_&�Q�X���w$�I*[b[gTB-�����7x#H#w<�C��+��i���IḚ�v|jM�����̢@���Eg�3gҖl�%1>��,���։�Bj��qN�}0�="z�KkO�]&�<�2�E߅�9}>��¨ZI:���i-�Q,h���c��^h4��fތ�1sY-��W��m��gyԲ�u_�����g��jBx�h��a��q���08�/� �Z���t]-uU�uj�@,����Ć���1��Ͻ��Ə�+���nS��=�,ٔ���5���w�.h������권�'�,���q���Q���ubg����~�0A6'7	ǌ2?��j�e�E�ou90����k�Fh?�9M#ʀ������_˄�XI*�����oS�M�tg另F��`�|Z��Z$r� Ω�Y�S��$TRI�K��C4����	.1b��^�a����Yô�`�׷�kAN�Mw����/ȾT���D����ӽ�}���$�D/��I/�}�����/�?����WH��1�L�Ɋ�e�Bn6௙U���%��/9���/��Q�Y��E+��!D�ɿ51Q߃9�ģ��茶�}[]&��HՆ���LC;����)��:��E)[
�ȥ枏3�4`��� ^S|�8ӏʷCle"Ӳ�v��0��hن�s~bƚMΉ�TC��)�lO�C�
��o)=|=k�@�e���^�ȷ���GMd��x������ۉyH��y}��DN-��tEI������SA�US�����Ǽ�>�9��SJ��D��2:]��wPY�_��i�lT�k�9
*��>LN�ܢft �WTw�I����]��,�.eW� ׀���]�~^��&�#�~~������_���-_��IXP��H�0��h�y��3���:8&0�m��8$S�L�&���?E-��ME�Q��$
I��6�2��$}���=q�92Փ?#����="���8����L�!�� =&J����%d>�L5���Q���㚜EUڙ��'w�9�P�����5
,���[�]�8���ֻ�g������r��� �s�Հ���@��j9+�c�t�>������M�N=���/�g���}������&�U�d���7'X�����̚;"�	���V=��#c%�&/���PN8�*9|��UOh;�b M���ġ��H4�` �y.��`W�zq��aF��wM��"��av:��fl��z�W�BlƂ�į�A3 w1y��b(�f@�6XkWZm|�{�2B=�N4��v�[߆̆[�ڒ�^��f�=�[�L���W��9g�qZ����Lc!�z�TU������Q���A��,�|�L�����s���s5�D*�t�}=�)=���j:(�lz�)��E��������]�RnY�[]���5|z�/���4�gJw��Et^w'n9�k��U�KWV&.�-���N�&[N�z#�N�<
��o{ܵG1k���"��3��o�D�{��K��4=?Zn�0�|��2��'�NĲ5Z���ױg��9���)��Òn��~����MVw>��.4�ul��j���9�2 �>i]o��g�\�/�x�ֈ�O��C��IAS׏'JI��bq߮�0��k�S 8j5���WMWPfk��dڧ���L�̰�V�Ӹ����j���� ��1���î���<1�t ��� TU.�r9ȝ�ǒ��@����2�j���M�����e���}�wbmQ�ț�&J I����hRqv��ź�Gƕ!BK��6�J�3�h���ލn
:>��@����H��UV�½H:L�X0��������R�J�Vpa������OJt��}�5�(�CF�����$�%3.�!˱����2���ƃ��>¨̵3tlbl����ҠJ?+貈>���t�d�_/\V�˦+^ץsl����Xw���Z� ���z/�!GRx��=�|���eh��EE?#���Чa��N�����$��6)afDH셣���Xُ���;�G����+s�l�x&O����<��:�5:��2i���*W'�%��4-��ZD�N�:�e�h�O�B�z��mp��Y����Z�4��?�a�v��6�W��@��o-��J�����h��3�h�s�1N�;��aӭ�R����$�΋�6�	T�K2�Ϥ��$f*s�=���Φ�ۅȰ�WG^ֆScĳ�,��.�~�4"&���ؒ�rB�M�6>"������1(�3�.%g)�s��7⹄J��&�6CMg��Ak7l`䨓�A`j���,J�y%��\zW�i�z"͡�B�H�@�d_�u[(�����o�ȩ��p�k(�|�RO+�"�b�?!���(�[V�HQ6�]4 �4��ůX:��r-g��'�D0ZZ��qK��t�8��0&�/m�r�D�N�2HQA���X�I�y����BW�;ĵ�0����hKՌ�CVG�z�+�����uA��-�p~Q@Y����x`�����1ة�8J�Z� xx��!̯D�첐����P��.l ^dog��1��wN�hNo:8

P_v��m��-˭��.u@+����(Ɨ�!;��9�d�'2�N�1L����G@g����SJ�@2�V������b�G+�204%v�M(|����G3-�6!7x�/)|b)bm���7�Bh��qv�VW+�3ת��ig������ʴ@j ��io�Z�59�i�Zh9L[&����0P8L���&0d
,��nY�w� �4h^I�����ɴ�u͉�}�$]#y �k?p���A*Ui�t���m��Ɍ!�U?`�z�g��쉶�ݼ�=>��j����|�˦ۧ�3Wީ��J�v��:��_-���S������b��E�l�s1�(Q�1�����]>��}��Eꀓ��P���I��&�a�@�\�5�|��R~��K�w�#*Y�1�[A����s-���L���ᓨ��1��L?~;4$�
�h�!@C�3���@T���%�t|���u��ݽ9/�O�w	R�w*v�P���y��v<#.ޛ���`_��>��f�7D���<	�3��Ct��n	k	5�r��0?k�h�y[�U:��!�2��ߦީd}��Hes�]w�RB�嶩K� ?BM�#�ĝI��@:q�Ǘ��
��	a�)�]�����{Ln��Ԓ<��1G���+�����A��!όb-[C�U��$���#����±"r�ٷv�	��7���Mø6��6[���aܺ�
la�ZL��<�P9�2"/���l$7T4�쫅A��~���B�����9�&���M=K�7�w�M���^V7��*s�=�@\J�]y-k��G����El�@
y�� $Z��ōk]��&��d��9~1r��p�ǇD���ԉ�jD������#`@�3�B���uɵ�ն��E]���5�C�����ӻ�����}��R=����k^�Щ��	������e���ȵ+t?�{�N=�G��T�œUjꠇ$jM�F��Dۻ+�|	?R]��h�o�o<�,�IY��C���R �Uǲ�}�^�Uy섒�Җ�� � �Ʀ�^�j�����F�㑏m׈�cلs��3�j���������z'&1�;ѹN�v{�cҥ����s�^��-	��)㈕rC�����kdK-�ۚ���}�GO\QMPZ�J��z�^/N����*��WP��|}J�z�l�gՠj�f�3����F��VLq|�cLC信��o	]k͒#�=Y]|i�3VI�6	�6kx.K�CO~���nv���KKnY~%�Ц ���6����#������շߥ���U��m�-�+�Nu���2��G��nZ��>���y����[RJ�Hw��@u�̙k%uEW�d��#i�3Kv��r;�n��O'�lN0\�H��D���]2��h��_��b�Y�W/�X�?�0�V�b��J��ck�d{�������i:�gr���I8e���|wr�C����	�)����j�#bM�:��sY�$F,�Ym��e-$D��F�L��I�t��[Z4����ϛ^'�u�"ʴ�2e����*�~�v��� �2A�0){����f������W�d�i �]��8�l��
6�^0l��
�G�<�D�!p�(.@��l�_�$Ȫ`*��e��
�`��"�㝒�>��|����>nQ�j�cA/و��DOx����?rQ:=�֒���g�a(W�x�H�73ITJ�����l7�=���⨏�ߥ�qOU�����zM9|�H�)L7�3Q�}���~�rkU`O0M�-H�ܟ{��fJ�ǲݾ+�
�r�Q�]G��T�4
V[x6�2�Q�Gz#��ע�Gڣi�c�3�w�2y|�g���x>$_�:�ꇗ������{�;�=�����{V빊q�/$<Ȥ���X��b��G�A����{~~�*���ڍeh0ҍ�Ǿ�gׅ#�$���k#��!_w �B�8��Cϋ����	.9Z�N���q�/a!'�*>�����[����V8��%HB�/�����v2�n��h�O6�okYI�l���dQ�c�Q�tGl�`�FC�W^�{�xT��%��8U�C`;�b�I�l�b��l����C�Y	�:g"�D�̫|v��F;�G!���X���퓂_����}.PLw�,�O �c��(�kN��m!�Sl����L�T&�42"<!5�3�jrgq��Î�H��dیN�<��I|�{���8�o?eh��)�D�I�!<-Q�_�j���Ą+R�"
��]�C�����]�O�����+�nDu��Xm;���B�C�P&8��Ċ�A�G�p���hb����Y��<`~~�����L��ai��N�X��}���x����&@s�Ԅ�XAm�H��=�M������~T����ȳ)��L���vWD�Hk�/Q�Jʮ&9覕J�����yr�m"$#1ʬ�Wt�I��NX}F\5��B�x�[��c��׮�H��.����?y
$��cD׫�k��le�Ak8w�����(����a�@Q�P�ޙ́���2�=�f�,��<,m�S��W�1�p��k�*f�	��!�=��t��P ��\/J��s��=�J�� �4>{m0=�
�q�C�@��gc�������{���+�2ԼX�����Jp�E�rp$�N���{1)��	t�<G�7���T�{G �j��o�K��^K�^\M�z�67���� �B'���
8��4��S]O�g������;�}+�G�x Xd1��|��	��ۀ��_n��R�xdP
�/�����b��Π��9��Kr���c?�YK���:v�Tv7_X���l�{��2OP+�Q��L`�ޭ#-�4M���1"F¯��+���9�=JOR�j��	��H��HD֚p��v�fQ^%�F�xꌶ޸رҪd���/+�c֏�>s�9�bxQI1��c�T����m�Pʫ(pM�G�4IU��wM�J1r�g�W ��`�o���7�54~X0��i����|���RP� ([��8�ݍl8_D�x�
�u����L}�[;��:;�'���6�"��۸&���iBrȏ��]KQ��[Έ��BOUO�.e�`*� ��z8�UA�������!����'Ed]�pd���z��m�+M���B�`t{� �D#2�x���ϛ{�Z��)��|)�������f�G(�,�FAQ=�џNbW���{���4�< ��r�T��sN0����9�c!��G��'��s�uN�}���թ'ƭ���FiT*պ��f��U����!��������Gx�kh�A��b8���5������7lgz ����� �Κ�`iO�#�1�b�C����L9��À9���7���Ț��������΋��qL���±�bω��5���jJ�z�6oG�Ƹ�Z��H�\�ǆZMd�dȿl���.�1�q�u�-CS��$+��v( �Jm�k�(�86��H*+J'�@�U���FC�GTr�6�R��>�<G���|��N� �{��k��rZ�ײv:{Pu--u�?��-�Y�у�+F� f����{&��
Ί6��l�q=X��R(�������OV��ْb�=|]�M�Z�2�9}�
irY�͞fX�a]6��
�,��"	����,h��d%
s�����������$]O�·�N/y�۳��π���Q�"5� �X�sN�BBY�2z���w��)�߂[5}@��)7ݪ�W֖�iҿu��劓������<�3o�	�B@�+b�E�޾^���b��y�;�
W�c���F�:�+`�uۥ�3�����yٖ����l&�)3ֻ���{$a;Bx��?k}�x���+��9v"b\�Y�N��7�Rozc6�j8�U��^�����}iӢ,M�Ś�Ϊ�3?#��V��2��d=ryL�I�Mg(�]S�K��`;�i�W���[J^��$»���^���<,��P�X��+mnA�8yhh	D<���W��}A
��@���vk 8x���8��/�^�y.$x��QB��9��f��w�b2�w�A:Y4+u�+�������ɂ'�9�ˀ��3�̽YmQؤPA��'�`��K	C׍]�Z�WXcQ|8�7���+�w�3ʓ7�c���бl����O�O�Ϝ��I8������@�L�\W�����l:%M��,�gf�|���,d�qI�[R���U�ZÝp��*���卪y3�B��ބa��O��ov'0���z(���I��[���8�:G���s����H2�:X����Yr���^em*|a��wc^-bv���B��Z��0�tu�w�n?bZ��;�B$���zđ��"�����?�쬬��I�3p�.h�W��`/,!?�_��-6�A��tf0%�<��I�����:��+�&B<</z�u Ai�k_����}�A8���ᓊ�pǑ�hn�$2Q�D� �îH�Ɇ[��ߚ�!�~�e`	��ɞdy��)��b (2.ǐн
hK�|���U��%,�<"@O4�zM��ɪ�sy���nB�=!���\^�e���&:�S��8��V�UG�����u�G��D	/�/�cg����lrѹ<Y��:�� H-_dOp�b)���;3r�0�|?K��X�����,��Múe��H��Y��[�aڎ���|��Q�o�	�����v�@Ӈ�j2����>�Vܗ@�踦@Ϳ��u|�K�g���qI2	^��&�)��lb�#$,���-� ��b�d������x	��jZI'gE0�U`���,��y�#	�,����Z��EcS��к����f�U��'�%�͂���q C�l�ȈV|�o��W�ԕ�kp����<����_^ū����p�%��w.��Y�*���:����_@�H�����bx�)a�����q�0��2	_gFد�[��A�؂��c���t+��j*-f4���|�d��b�Ơ���|6��]�.�J7��њʞ��]�!27VP������l�U1�2�j/��!�c�t\�7J�J�n&�;�֘�R�W{Í^X`X���@�M���=�x���l��*-jG����2�+��d!|:noB�����إC?��;�L2�.	�yT�J2�f~G��:C��yae����t���2��.��Sz�3�}��~]f�J��p8Eg�{���� �J�dnr�Hw�	���X I�dII�>	��V��pv�O�ʠ�HB���{�����ğ׃��MO[z#���">��?ʥtg3OGo-���_�Yɐ��&�`�C��*k��ߙêO���fՍZL����0�ً����$kTuѰ4�vj�4/��D��*ܷ�f��u�����{JOsYm�7�N��s����TeXD����� �=;ٸU��I��l��T����+�Ǚ)yl)L:.����ě����j����p�%˛W��[�Sp���+W>O�����X���qe#ܺ��L��D��+}�I���6]��A+.C6��ݖ��DO��m�J�nE�Aq��+l��$`C�^p^�.�:�mr,��o����3�$��pl��I��TgmV�|�qH܂ ����O+~��0V��=���n�l�M��R8����o�v�Waq`o�X�<�v�	��%�j��#���	{�nvs��`!��U��2��{2�XD���� p1mSc������z,2n.�i�wh7혬$J�,ʠ�q�&�����g�tI��dV�%�����iꩽ���$�8�Z���.ҝ�Rl���/���Ϯ5;R��1�sGu�_�0�&U0�ŠW.*)���n��s}Vߗ�"y�� �xu���Rc�"���tCZ����~�~��)כ�5(mP��w��]E�5F�Z�.���s��M�Gb!��Q��܆Z�l)a&_*6����F�+��8�����r�qc�����[$��^�af��}�����h��!t��3d�V�g,�ϫ{���օ��_YT�k�s�'��~��҆#�C��]���t(�C�`-����+0�:�X% 	�<n�kF:�n��+v+qR"�&Y�D_��7�g��	x:�g�[@�Y���do��=�۷W��>`쭴0ҹ}+�Δ�z,(/8&X$�H�}��@.�I7Xjڡ�x��dk]���*Sw$�Ay���gu�8��tiHK�(GT�wq�sAg�4�߫8*��(�0쪾��cA��Q���i��M����"j7Q�޺pa*f�
ɖ�oU��=��[:�<�?�[䍂["��>*���\I l�}���.#d���W�{�谙��C�#l��r!:�CP��B��v�G $���͐| l~��1��������l�CD���{�r�U�@�= ��9p������C\����7�*�ƙ��I�!�r L��J�׍�g�Z�w.`��%�Yt}L��y����Z2�~���=��wCw}��!��\�%B��MV�)�+��2�>���7�K�	�j������\�JV�}/U�w[��i�`���pw�fo�;�ja���gk��+��!2�&8I�O��6E�bbӝ.$��qrE�ȥ��T8�˟�Z��D�p2�)��ke��~�_�D���ĳ�_�:@��+p��	іIk[�.T�a(�������	y�=�8k�A۷�1��4�N[^�몼�f���H}����ϩ�|�:���(@M�	+�g!28�V7�捬X"$�������렰�Y�؉���Ti�2V���<q7��w��k��pY�PS��(t�bi��'���@6�ظ=���\XI����`HDU���˸�
�3��+�SG�dV��J�>�,$�^�i���a�Y�(#7m�#�ؿl��{|B�$������A��_&����s\S�7�pp���<R\�QX����?D!��x\=�K�<�q9�2F�sCnqK�����}���Ʃ:��)����1�E&����x���0x��!{����Aa�b����.�>�d�/��"g(e�-�%�[�W,���lh+ �yp�����E�;��~��O�;f�A�����9:ۗĮxH�W�VD������Fæ�n�`Y��B��f�}��Ć�I�65��7ה�N��(Bk\]��"gׯJ@�a��ţ�"쌻�:^�eO]�Q�`n�0�R���re4)F�}C�7d�Q�q����f��ܾ҄����yl&�wD�T��שf �R����JĨ�Q~�ݭ����	'�0kyb%�Y���{Yۗ��{7�%�k!.B[{��MY����3�*gͅL�ƪɃ|��2��p7B��eIs~W�f	i	����T�I�-�\ui�^�wH�OT�0�6��M.f�Y)ұ�.�)��p�����#� z�l!�J�pF�cs/���=�o�W����v�ii�*���Cf���jlz�k�*��Ӽ� (�"L�c�� �c&?3a��ms���� 3��;����xq3��9()�gJ�����44�C�a�2����M���v�$ݔ��!A���,YQZZ�R�?aJ�,�*�' d�����"�h݆S�T��n
�����G$.����`7I'[���́��0Gq��weR������Y�W�%�C�[�]K[X��ڋ)q�Ǫ��MP�����k6��ʝ �eL��y����ϔR�y�a=ݘJ� ��U�0�1ew0��C�!�f�����Ɓi�I�^�H*�F3��X9�~䬶Y�g�ҙ6��b�ի��C���R��0t	�a�3�s���؝����n�8-�}T�?����(W)�?S�0��#��RVx^[%5�9�:oܹ^gad�ޚl2l�eQ%ľX�9��.��Z���[��߀>�lP���:��� 0�G��?o(�|A�XzQ�9\�a�ҕ�]����m�X�;�
�l���CQ3�H�-H~�@b<44~���!>2	��)�NM͞y���;� 1nD�ś��-o	����F�ojUtj=�Tb�yGR�k�\�AG6=�r�?���X<�hڤ���[�b��9 ��`]k�WT��e��&M�٠�,$'��?}�$8!,�vŇx�JԦ����
�� (�wӺ�]���-~�� �9,�R.�Mq���F�����r��H��l4>��R~3ܥ�r�;�MP���X�K��\��������1���6�.:�N�[]һG��|bFS\v�T�k�U��P�:�OgT��H�y�"��l�ko�5٤���@1�%&��׉�L�a�Hi�4{��C��u�a츕�ۓn�{�P��L�<���>���PF�o	�������k��k�߅�[�b���i�ʅ*�>\#�w.�׹�sT+���ZR��V#i�n��@�{b$:�q�#\ݍj	ֵ����[3r��D�g���\�8�r�u-�k�+����>�=+Is۹A��7��Ii[(L߽�嵪F~��a���Z
�N�]>�͈��&�(���U4�磮�4�`W<�C����"4��:~�gJ��O0g��S�>�{�G��ci���|HqS��Z�C�|�"��z�l���îavx�.d����ϥ�����Xj-��LK��/�&5"-��"?&Hsa΁��%�j��߷�q�l�;�-����f��yp��t�F����k���Sh	-,Va#�knT�,TFVT`����0�2�T��f�	��b�Q�E[a	Z;�����������R1Ͻ
Gj��Kj"_�n�q�&������a�sݾ�t6/bq��ɕ֨0�r\�-E� �5�^i�����*Ȁz��B45�,��(_-���u����b�����@ޗG�K�:X\�|[Ƌ[�Ȋ4�.���v�B�G�Y̴�氤uA�
pg����V�K�� j��P.���;��S3¦���mS���<m#�/n����a���t���!���غ(�{f�܆��aJS�0�r�r����:� �Q�w���6�6F�'](-�����h@���wk���'��a��-v�vY�*�Af���y����͊��=�\��W�(��f�� &޹�%��Gۧe<o��P�v��|z3�@[�l�n����@����v/�N�L9�W���Ű�_6���{a�*�
����(��N������LDY>iNġ�_8�z	������B%�y��@Z@�����?#���-(ٝ�i��I�]�VB����̓��Z���JX��d��þ\��*b�< Y��¡�W7B1	!i���j�����x$}�D�ɀ*ۦ�t��/(��
�����9X�<�CyF�?37�I��]������߷:.�ȗ���d�DASzW�Lo�B��J2�S0��,���K\1m���	N /b:���]D;}���U}�~R��#W����s?�o
������˱��Nd���l�B�!�JM���T���U��XAA��!�16����"f��n����;&"�#X��<t��@������'���UÍF=u.(�GE�OeK6��$��U�\`���ꐻ�7�D�lj3�=T��4�GƱ�'�EVu��������༇a��k�y�^���*RP��OjRX��&��$ߛ&=���/Ȯ��k9�ч3f=�P�L¯t5L����L�!"���M�+��;W ����a��p!���W��O������� �Y���@��6���>��q�20D��O�"��{�)��\5����a{��i�d7}���?��^gݽer�z��8�,�I�^�Z;�����@�L�Qi�9"��8dt��"�A�B5�4gw8����N��xq��e����F�h��A�'�<���M�/�蠪|��H
5��-�%�V��,\3���<Sݲ�}d;<*�@���NCz�wO��KG��o��>�:��[}�#���n��S�'�s�8��t 1x{��N#^Fۋщ.�Ԁe�蕲���u�������'�Ёj�ю]}�2�y�3�������Z�7oE̗��<���Qz����\ǘRR��OqzA�� 2|�vK���g�P��nw$��ۈ3���q��,Ę�R��e��UH�t�e޴�DX�	���YIh��E�d���o�O���M�Jm��y&�9�Y�:��a�:.��ao�a6�2)����=�����6�
�Y�̉lm�/�h�x���s>����|	u�m�/��S���F��TB^$Z�PAyo�*�q?��U��|��!��^���2w��0��I©�3<G����r1�����������E���rChM!�B��
YeǦ�,�A�&'���tCN�����S|Y���S���^�3߯R:=���!7��aό�q3ӜA���y�XY�:��,5�no8�l��X{�p�K,G�3��|Wx��\"X����"����Ѳ�jo�llD�tW�ܽ'���/���!{��T-��5E�����֫�˖����XN���<�;k�h��!T�A\ 3M�H�#?�Q�ƾ��m˖R{p�O_�(0C�C���#�����ą�E~�2�$��?
"�8�u�֦}�J�-y�j�D���?,ȬH��#Ç�Ɓ�c65�9���O��.t>W� &�BY����>���<O�G+ɚC*	s2��K���e�%0�!!�"�/�1�?@9�̔/����|W9��o]6�u��ZK�%�t+�5�Qu�a����F�)g��?<'�0�+�~覿�I�Ÿ-�-&�I�s4���Ah�f�*�J�*��;����"F��£�E�	F~E�l0+���C� @���������v���߁*���ȴ�Ӄ�nTv���_��62s}`PXO;l�̘�FGzB���\���ěF6M��쨼��I1���\Q�Ԥ(��i&�t?o?��ξ��jXI�<	��Q~I�+oF�UC*��ȓ��=#�7ϔc�}���D>����1���e���Pv��Qs���N[��3��M � ���5�_W?.��J{�Ȗ}��"�~��]>�R���nOm	�A����.-0f2�1���᳛Q?N���*eq�`�eE���t��r���<GY�]�-}H,vL1��4��J�G�
��+Ȝ�AE����j����)a�2qRe|_��޳�0*M�,�0�E;�aq�n&���_e�C���l�y�.��[W1�YR�H�9ʴNi'����t(�i�������b)0W_�F���Q�,:mrJ�z?|R����;�ڈ�V�j��[��Pv���Xm�Sr(�[�J�ee*���>z|�W$���Tkh��g��r�%��L�Ԍ�B����$�k �PX�������y�"�sg������^�fI�+�L�P�&�I��Q�����X�����S;���%(���*�6<) ��Ӵ:�z��C�6	6A�u88V���K,���T�D�1ѥ(��K�4V�V�B�,��S�O���?���D����:]�%��n��Z(J뙡c��4|.���Z\��:ɚ�z��X�1�3Zy*l5Z�T������1�#�9b�_L�dMN�3��z���@�g�?�y��-����o�^�O62�t�&�	��̠@��>�jl$�fgL>�]��u�cҋh|
�=���C��̿����Iqu��V���~e������g�D&q\Nޟ&&Ə D�m�(�'p*¾�x�X�b�C6��=Ue��}����HZ�T�u��{�Dw_%�^L{1ؚƾ�'�,�N���E��ة�(	��W�}'��ܑl8�l���sq�������5DѰ�����r,�Կ���b�i���o~k��3��}Ȑ�����e+��u�c�	��ki^���".zV��p�:�M_�|�ů����>|���"��҆�h�sF� ?�nW�\+�o)������h�ւ:]�`�=��zJ�Pk��ЧA��]=��&�4y}Po� �=z�)�z��G ĶH?�#�J�}\{K:"T�J۰U���>cC��Y�$��<���b:�',�&�d/���߾~��c7A��5�`;h�Ɇ��Lf�*N����j>���]��h�7��r��TP�M8J���Cl�Pd~'��UIi�rG�k[+J$Hmzh�A��aD��y��?�&K#4��9<������̗u�y�����K"����~�JB����,9ۆ�:-���hI��<ot˗��~���9/����1'�ap��n��}}���������\���G���۱S���zߝ��o����6��i���Z�^t�̸;5��w��aa����O��Z~@�Ƚ�����	t;闒�~��@}�1��
�d�c��Э6���PS��G���( �c3.CΉ��������:kp��/�T�MA�P�͙��lQ��/en	v&> ��љ�(��1�Ԍ��!�9�M���0�E`���H(�lj����ƚ���OT+lewyA K�`�؝n]pS�ҵ���T��D�)�/��kaOz�����cB���k�U_�7O�W/Y�\t�kl�HkE�2݅����=�ܷ�ؔ�RS��Ai��N����x	��<�p@���9��숳�kDPj��BT�����2E���<^�u��B�IҧF
|�Z`��x����g�"�4q]AC�k�Q����l��o��F�C7غH��4�b��|�.���ͦ~}�H�s8���>s�8�f@�k��=����:Tk���a�k�b��
V�ł ��7�?��{ϯ`p����Hw�a2e5 @봾a��6�2�P�ݽۨ�|���$�(4��W	�##�wW\A~�*�6E#W Y����k$�A�q1ax���[%2��	�^��1��g�6&�!Բ���6��?6��a��un��_�ƱМ��@ ��ʊa=w~����-�.��tg�sc���]%m�( ���C� �t���St���S��w��߀��ךH�l.���� �T&��  �|g�\%�)��Sگy��f�$�Yt�o��1&�/_q�{��woBށ�(�MR>ݑ|\�;�]<������tܑ�*��+�HD'Q44�Q0��s��/����k���mu����'����!Q����TX���P�;�i㚰	�0X��AK�\Bi�^���� {����Q�6P����~�ߗsua/��C��Q;�ɇ�.u�b�]m��jz��m�\5M�����?f`^8��[²ĝ:��K��Dq�A&A0yEb �����h�^�ڐ�|�e>3_�23l4��>PՂ|�*��������u�M{[=��Dʾǉ��qnP<��n8�h`����ɟh��5pO�%@W��O���6f'N�����V$w8�k}��1�e���+��`�������!L��NGY�+q� _�Q��'���C��Fw����;hIv��^Ր����=뱭[8V�Y�5p�Q[Kx�)^���KEL]ƅG�O""5/���	�"=�:YtA�<��.�?�,2��qØH�ypFV�-�>OT���L�\{{��fh�F�?Q!���t&��A�ovo$�r��'�2.�����LU�LÔ+�{��!�dۄ븕�~kp���2��� j�7���'/k����G�s�����G�+)���q�n�k���p	�B�Í���2�&�	t.����x�N��n >�*�a�9�l�Z��2�:~,�a�]�{�$p�6a���b`�*[��y��� �Pi�d���s�@e��̵�x�&&�������$o@
�
�/-���;���ې)���J�<�m�H��vY�
hAu��%�^>�R�o)h�7��X�j_�g�����16�W��"'��k�5;�@U�`�k9��J���W6NT�n���@�Z�~�MT��U���s�?�Pz�����Z�h�� $OϜ���:G�op��DUϭ�?EW?"_f����$�徊u�k'Ԇ�z�5�A��8����P�,��a�4+(C������R8�Q��;�k�ik�$�0|^�Uiq��i��~y	��&��Di�O��I �����"���bƉu���쀭0>�.U�Nn�r&������
��NPf�R���!��^�_K�|]�<����fm��p��?�I�h����,.!i7t��LW��y�{� �E߮���X�s/��\�D:�&j+dޫ�d����Ɩ:ZcG�.��/��&oc��I6�i0��\�C>Mow�B.��
)�tb|��]�o&K���F���w��7�A�[Ʒ�d���<�u�"�u�b����^����� �����=p��0�*r��4�$z.U�V�@��1��'*�.�4���B�ʆp��G��#Լ#Qvb+{$}�!�FL&���`�&�F��H��)o�~�.��^�B8|�So W�R:��4�E�1ň��;��E��y��gk���B���6�u�9%	�` �ܴ�d�#7EH��<��ſYaJރ:F�� $y<ס�_}���S�\t�]���X���9����F��rd9�tv7>D����Ң�Xgt��0���5��n�@=�Z_���$�ï��� �.:�m�{�K��(֢��|%ۚ���0+�j�}��|4�SG;����	o!�V�Rg�B�*���F`CA,/��� 9�s��Q����7&���ctRtnΥ���"�<(<CIs�;��\��,�=p����A�ذ(3]WXVҾ�V�� �9��!ȷ���K��I<�U�����N��(�a�n��i~X�qIVWUB��5�H@H�]���p}���n��m�M53�$2�	�w��� �D���oV-G��n~J#��}�'H��d�,�q�
��tx���H��B,H)��Wrzq�@�B��X^�= 9��?��� ��a�"h��,{%��qrT5-^}�9��l��+����J�Р�`�@�P5�ƭ �M�z��e�m]_�ǨT)�J��y�O�P�>�xHߕ���6��m��n*Ԗ�ƕ�� '�E��C����XD#�|�	���Gk친�h�����)u�"��b߄��� S\�[ ���C.mr�u�b��2�p�[uN $���Xk��wb�ķf\E5�+��R[��)���V� *0< ��<V%24�T���U�����$�@�� E�}�ȇ��c�_�����[.^��:ŵ0���ҝ�nu}��>���U��m� ��+o��A�V0����0%Et���kny�����- pE�K[az�9��zb�ʴ�p�>V`�����:xO+���$�j�w�'�#��\��x�]�P���jޒi������1��/�J�n�����s%-7��@�{K"S:�L�2�@R�W-�z�j����{Ȝ�^z{z�E�(�)�/�"σ���*�|�x����~��r���������T��/�� �G>�A�<��~)��>�m�>��`Q�)(�Pr���;�����ѡ9}�c���EhlaJfQɚ%{�L���e��� �x-�H4xܲ����r�|�Y��4�1�7�����c2�����>�Ǐ���,8����g~����Wޘ-'�`d~M�T�oE/����l���S���X�,����tܾI��m�����`F^3��&�/�}����`g�vH�5%���m`��x��K�a��l����s���C�-��u�Q�V����,�ĳ�qy	��9�O�Y7�g�~F��'�4�~%���U�Q�	�o�H��dg�0��.���/Y?���"_Ql��@w�2�z�G`�o���SsXvjJ(r���0�5%���#@q;�X~���i �4� �LU.2�eIĉ��.����>P����,H��c������8ӎu6윿3�H����Nc9��7u�yr	ɗ?K���ǟ,<3͘� ?�;q�ϭI�s���y~�����7���b�#/N��)-�dl[e:���cV�k�cM�����ӱ>"l4W$Bo����_��ϭ��!�Xw�P���,}�Up���;���H�C����!h߸��l�m�We�D[xyP	�ܰ�o�g���,�;F�q���� A/k�/��-�,�p˞"1�M�/�7�=�<I�`C��ސ�TGu Ҥ����gQ�[�Ȃ�J��`�dn־g�[���c�^�M.Y�w����2��H����m�!�A�婵�	�]�)�V�O�e��d��qO�A�x����^���'�7V+N1N���g�%m���������P�_�>	����Q8�7FN#S�Qq����u�x�&��X���*��M>�;�������_�$>��Xjj+ �Ħ9�@=�DF�?�F<�g!�P��?����m�����I�,��ʔ�d�/�|��מ��ݿ�9
��_Y�c��/�L8m��%L�5�1d;t
��P�/>{h)�Z���{���H�0
g�%#��)��/���Y����-sv/�+S˄��UU�M��F2�Z�M$�.'�/�\���o<|��kǤ���r7u�2���v��1-���G��8��Ӝ��x�1�p��+h�{�<v���F�#!Z$z��Q�=��_��t����!�S�+�'���r^h����C}�����.�w����:��p�c� kJ�6gs�[���ox�ٸ3��G#*�/ؙ8P�K;�=1N����ި,ω�)�U�Cq��q4
�r�"p��A�Pc����8*���u��>zh�1n��g���Ns�t&h��@�����E:�$����;�D� J���v*t��oX��>Vƒq?8Bۑ��h����g��ԕ���_�-�^�HJo4�\�)�>�\>���KDMK��[�/����;� %�ƽ�&��A��.�H�8��a���uU�􄀴�a6'W���xw�r׺��JP�s�KI#��Q]�5O�f���|��q�RW��߸.�P2O���t�LM��j�?�H�W���3���jU2k��&ao9��qB�ß���������l��[�4���a�f/4L��;b_���iux��ڌ�qw�P�l0���|�Wœ[��O�ԃ��^|;��ҼfP0[��$��ڪ�R�^ դ�bo��f-)8�Nl>�Afb	?O,u�N�?Ge3��[�%�@�����;>Nz �45�_���P��I.V��'��Q���u��/k__�WoL;�t<А`�F���K+���1�:���L ���mp�(;�Q�v�E&�4�*p`h�c��I
vyb�W->���ʃ_�XfX�C�#��JDySk�$��X:P�wd�<)wF��d��h�@�]^K�3<pۄ�@3z�6f��)�8i�z�	�kx��q2]�9o�� ��~WD-ڏe{i��Ȇ*��	mW���SU�@�G���p|����p)�̱x�i�.;����8�yY�dg�N�������ծ�,p��lj�Oјҵ�-���f�%CWt�)�y޹�\e��u<��͈Np۽�*�~�!�ΘrMʟRI���BOr���k���&ܱ:
�,pNxb�z7po	+���5o^�@Y ��Th��F0 ���0T�*����T���\����Lҡ��5iF <�h3�/}p	��0��;�7���D� 5ܤ�b��fT�e��,�Nc=a���.v��<o�g�m�GxR��p_���;C�(���F�Q�Փޭ�_
e���������b��~�{ԟ�3of��(M��H����L9�͚w�""��>��:�Pd͖~L)�Y��υaR�!SL�ib�
�w�3G���U�=v坄dj�����tΖx�w���뽺�����{mJ�b�ijl*�Nd�S��U��1�TV�KPb+�۞�N.����P'q��.�~pР�f5� U�V���d���N�ٙ�����X�mF1H��%��Όt�&ӹ	���d�]�X_E.܄s}9g^�
K�����0����R1����_<7O�T��Qox�Tᦝ"�/�+6C��9?�K�9�Ȝ,�#:;k����J�}�w�P�>�;���K�
�<�wM�ަ���LS�����
�g������'cR���k��=pb�G� So��Wn������V}�Y �&���Ú����Xg��,��]���d'*�y7�zE����{U�,W�\RM	�-.:��q��؞^�F�j@�f9zZ}�<��ua��Mng3^#l��Fك����{���E��]qH����Z�c�����N�]�Y���=�[$��&&V��0h	��>�B!�����!B�	by�{/E�S�ة����*jm}a���}�Ċ�bq��8��[����>�<�w�Z�[��.��;!�<1�免*��,��������0��鞀��׬��c�8^ h�c����N��
6�/��nC	хtw��`W1� ��5|/��Z}]uQ���;���� ���F���-�oJ�g�p�K�K=��đ���l���g^�C�z��{w��#�Ǡ��Z��YHa6������m�-1��M�	,�Y�d��"BB�.����=y{f-:��<���$��P�EYbl�7mv��FȹLڙ�i=�&&U�~���[��km?�9%��˦ʿ�F���ӫ�X��7%\�ҹ���	~�Iٯ�y�0|B��[�Y���d�؉��)1o ��Q�I�e&��h�:�c7�$�3He��Cݜ6�zu%�h ��z
���zS�]���%Co-�a��m��DB���`G�{���
��O��>�� 1�UV6�|����:Xs�vuM
"��a/�����5�����S�@s(L>��O���>�L�2ˀeO��YՎN�c���o��J�V"��T�؄�� �BSL��?��
�A&=S���n�Ě��T�ͦhFP5ƻ�y�����6/WE+����hlB��Ed+�(��+�'q���`}4<jR� �����1iS��n�s�����@�]�4q���\�t�Y5u����!�k����rg��:M�tiSa�s׾'�Y��h�|���=���]a�Vz������E�G��=�rj'
���lU���1�f�BB�7�D]���DB#cmE���q����МO35;�*{!-�T�g�tt�j1����AE�qM8�0u�j:)t���Sj��1	+x�j�	?A��\��P)�\g(�v7q=>n��\��U]���i,fp�|k�*IUƔ�J:�0�>2Xk��)��xDX�o`�恵�(Z�z��#�Ey9}O����i#NR�Z�%�,<k""�[�wģ��Lļ��-�6�w3[t�R��2�Θ]�|K��Z�#����&e��QPW6�YAL|�!��Ř��[}oԦ��;^�pP﨧&צ�C)2��
D�6>��=�\����`�	X���z����9�!\�ZV�Q|:���<+Tω�
e,A&*9B��sPĹ��V'[B����|��(5�{�ʳ��c���PJ�W
	F,�4����ߤ��wb���m0��B	�W�:��c:��I�=���El��#�/ؿj�I�M�����C��."�U���,���
1���1D^l�U�tW�3��x�ұY>oM/������H'"˂�xH�fޅ�ï���o6�Ay�u�|gl	V{l��b7�����B��� uC!���/*��ub8��.��I/4!���D�K�+Q����脇���3��4���J�wn���,"�P]t����A�B^���%�ʳL%j���HN�� M!�Zr�c��QH��?�{�C=݀�HA�E{�6�o{���c�#'�����rAox|*8���]Ȟ᲎�9z����ƾ��vA�~���e��Q�f�ȴ=�J��������0����Ճ�Ό�o�kd�7��X�G�Σ�q���'������v���߮���]�B�]�Dۆ�5(tW׬�٦�PU�S����g~��6�w=|3�#;4�D�����2j�S\�3�:����j���3s'�3�ln�*��۾G|T_��[��p�~5�
��IH� ps��f�|TxƟ9��>#��ɡU?ȶ
��}�"�������$3��$o0 =w/��J_<�����냯s���:�' +q��4�P�mu�h��w���x�V_�7���0u�$��e""L3��i�f@�M�ʾ�z�'s?8T4��l?��/�Ĥ�"Nt����e�08i��ԋ�t�E3Ҩ2�Q��� _�V9C�}��X���'T����SB>����L��0��r�c�Q��6�- L�lV��6�=���n\�N��3U���%�Q�#}�Η�T���F6S ��!�\%�c��tf��P�Xo�_�0��״�"��@"�wf`��d}��R��>,)]_�Y^�Xj�W�I�>m<
�2:�؅&�fTQ�vƩzJ�ym_��7��8�qp�4�]�2�w'�܁��
њ���yf��I�����Q��A�	� %=���1�<�욤|�[�S�|�zWhw�Ōt�rG.!;��Q*(�K��e$��\d0�sT��A��/�h�w�u��v����p��ߙ4��d�w���Ђ�H��y�d����%��*)l�鍟	�:ڪ����9H�Q�B�r<�D���..��+uRJ��p�7!GVK�&U��E���oEJ���Z��@�o,��H!N�w;�|���Ų����8��!�@B���5:.PB�1� ,�GZ/php,K�ц�	�><3t7d�\�:�}�dW�N4H9�0�>C�������)[�M�0����mU!��,���EL�S÷xi��/*�;�����KB���k�Q���Ό!�[��H�m�2��A�f��5Jj}~����m0�LWOfg\�I*�Z�a�Ƃ,eiz(�;t
n�a���
�.�����&��,so��5�5I+Zfԩ���b
���96f���\�(!�8�I�^��vx���(�U�J'�,Z��ߛt��)HEXP��M���&"�Cܢ�C7LL�]eD{�o�5��S��,`">d� ��v��~#o--%0�Ӭ�2W����S�%����n��$����ECUߋ�&/��Q�?��>Ms�$Z2���T�$�+�P\�+Z"!�h�h��ψ�,#YL�B�*�ㆡ��~cîU���5�S4���$k�MFh��b�6����Q�^�$�"r���}��s��T]��0�׎����_��Y��I*��-��Z{�G�Jl�[71G4)xI����A�:S��а�1�����Pnݑ��A�9'W�t@jƗC&V8~+d8ŉ�]Y�0�8!W5�:L]V�m�U��Z���=���֝�������KP-�h�L�X��'�y���\v^>�`��<�,�ћ;���'�e/�-��ǳv#�$��A�"��[�{�|ФeF]u�:9�`3X����7t����ee����#�5���K��sν�"Jl����@Om��w�&�
�6��V��e[5!��]2�vAmf��Դ{����{������� ��}���BOz�'�3�Z5V�G� [��@ژeI��`��Cqs�ns�"㨳�<���4��6��ɨ�7�/1�54k�[�;9��6N��%��΅�����r�=���'�F��rθ6�6�L�X[�޿�a�J���~O-��5\N���N5B�
	��G�ygy�^NG�YDe�a���o��%��dX�B�V�mm1�Cz�X�~���4.
�{ \�h���?[�X!�͹�f��^�qX:�:��1d �*��p��q�e ��
�)�",��A��j��u���	ɏ�ɜt��u]j��U�����fG�xA��
�}�����Tշ�{��{?+��w���x�x�9J���p1�����7Ӥ}��"Û�����1Z�]Uh�m��ɵُ�@�6�ǯh�+��(
s���,��8z�x�e���k�����)�IoK���-��V��s)�!�q�2�+ğZ���;�aE`&
ˢ�����k�J�\�:fA�t�1(��18�b��m�zX����o~����F5-���HD��B�(ു����Y��٫���&�;�j)I}�(,o�E�t��1��
����9�c�¤��}�L+s6q�Ghv6D���˗MTx���ǈ�����X����GX������{��ȞtZ�t���F���m��\�ctzO�2hT|���Y~=�t4���Ԁ��j����!PQ����l3�C@{�M&F�	G��)�Y\qZ&�����c�/�g�^��A�W����M0� �
U<Fx�6�r��O	�� �W)e����M�;���r~j<X.5x�ַ�s<�W.� �n[�Ğ�q2x��t��[o�%̀�P�µ+#�%�'��]L<�狼������ϝ-�r_��#������#���p.��ŌK��l�ew@���L�_(�^#�����*��\:��2�5~�����ƕ��郦ݫY�$�%i�vs��ހ,]�-�tU����Y���L���le	�mA���^��X���$a��1�z�nEL��zc���^d6F�ه}�O]vk亴`��X�]�2��X;��łT{0(�9�����d�[��o������	��_i����r3�&!7I��[C�-�_6Ꚁ|o�x���	�f�����#D�9-�^�}�D�N�V�4�;� Z���bh9>?���L��̤h�bD^#�2�G�D�W {��4Lߥ�=�[����;dA�?�ä́ȏ�����@�LYw��/�:Qsя���Yk�#���bG-q~�@����',�>��%���Di�!��4�.�xp�U*
6��0Ҟ�cͽ��;�%�B��y�g�2�@�qe�{�X��"���0���c�J:4m/D��㊧���f�����F���^��e����th��B @�;Ōnn�*�E5]Y% ��>�� �.=���p%ep$�]��������f�<�����r��=�ܑ,nX@�L�rAydN�����xm8��*��n\xV
[�k��'��H�>U��/Ӻ:����4��-}*!ɓ[�S�4w����������$]Q�4Q^:牵,y-I�7�欌m�J!����{'~MbbeM<����H*�t�,j���������k5p^�������d���b�j#��ܹG�$��2��媄��u��dϭ��9n��sN�#�T���{c�L)2�J��(�	4�HaBAC�*�}d�i���0#&�V,'�eH���g.�Ip'��+�����u��k��$lɹ�M�x'� >%�7��.N�~�9w���SO�~��q��m��\�S��em���I\�A�fu�8�u�@.��N��Y�Nlo�8/A�(�y4_"��ýX� ܛ`��k�k}��oZg:˸��Xr�[�a�o
��ř�YY�����Mg.���m����ֳZ���q�`�̺X�P� $o`|ksc6F�5���R-�� O�Fd�]QYY�$���i��L���:kR�h����}'	�	��\��&WD��L�HK�kl�06RZ��HB���Գ�>w�BK�#�	�*�I4T]�a Q�����h�ݘN=�E��	 ��y�O��y���Q�Vo(Ѕ�6	-��U��I���:��j;�L�s� (���aV#$���#kc오�n�PU����@�è���b��H�޼��������ɱ����%ɹ��U֗r�F�Z}��]���6 ����f��ٯ��Y���Z:HY6�!����͢ '$�#͵.��6p���azۏ�e�����P��v�r��IRwV���y3��3$6� ��������^�X��G�֮e��D��@m�@c��;���-87e�I�(�M[�q�È^�5(�/�i^-ȏs=6e��%_�Ӱr�π����dpe�g<N��y�?m}ޮV�x����`�v�n�������L�M��YE$�M���r*��pZ�EBx+;�;�s�=J' �ܯA��g�ܭ"�e�J�N��نV�_d�K�1fgƘ-YPt(��������J�s}��|ǩ��C�ٱ���{���kݲ���K�	�I��etg��D{�/��|�д`����A����k�rp��&��?Jh0�v�n�N��J��*fF`K���N 
ܳ�du?+��3���׻�����q�4�����薊H{^�$=A~X�1O�1Ӹ�b���|��I7߯�Ыx�h`�'��sD�~���	z�����CŦ���~s�q�ͭl���j$���vHx9����0P��l����^o���LƩ~�Ѿ�~9���j���I�-l�6�2.����0����{����R
%�\���,Q���A�ϻE��0^bz:��빌5`����� �L�3�r����$������<�ڲ3F�v�c��Y&��G�JD��D��S���.���d��N�K��yfZ�ʞ���׏��P/����!"l��WÑ��d�na#CZ��S��- ��L�^��Ô%�̀E(�/�����E�U�|���x:#��ӄ�d�t��̕-xɂ�D�^{�{�}�W�k�1�[4
CwUp�=���u7��a��WR�D�,�ue��Xs[��^p0�Z
�s
����C��6�d���;!�S��f4��&RnhjO�g�f-������G`q�i���\�1�{�1��J4�p����=�Ê{�i!��ň�^�-3�,�@ ��C3�MS�a��<L�n6�n�F2����zYh�pm���qL�%'?W����,�g0�n�[��v7�i�dŴ�K� p>a��̉�7�X�!�����(J�Z��SK�B�X�QZO&�
B-��
