��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���!<So���2��E�!�7���feI�R�34�F�\1uR�XO.P㤳��"����(W�����Y�LXN>#���[���٭{쉉�J�l0�s�ý�]ceW)*�k2���hj�i��I�&7�׀J�Oj�A�y&q��Mp�|���11Q7�3��+��t�`^�v{���.�����=*�I�6T�V�?��H�C�0�_�ҍwY�V �:�Ca)Y�x�G���C�������O�e�+:�W�5���Z�%��l�v�=m�lPZ#!��z���L��đ:Eg�-��9�aw=�R��ݤ��v��,u�N��o�'�oȌ���[����̬<��@�m��v�5OX)�,W���*� Pj9�=���=�y{78'���-R��H��U���uFݬ�6���*ֺ�dCNֈ	�8]2�8q��2�Y/�;ߛT2�|��B��]�zg���ge���-:^�O�x��S�2�����|�W>!�(�?c��QR(Xm�Uk17d�6q��;9��F��R֠����g3�㵳�%�q ��Q�oΛ�����֜};��	��-=ڝ�*���ю����|��7cw�:	ZO������_(��L�\;�>�.Ӊ������S2_���g͖��qh�%�;'���e�ى�Y�7�x��2byiV�Biᑸ!br���Pe�����n��-i��̜-�a�BI�,q(�o�����r�PdN(�n�@
����hM�~h�wR�S�AׅK	3I��T��-Ø�v/;���^PX!k%�0/6?N���H��ng�t�����<�B��8�%~��@�3�D]~!8�Yo��>�]����'T����u��N�I�f��gS�Ǎ�N�y�}��<����pL���蒼fm�x��:]~/m:1o�B+�X!U��!Mej�͋/�a�7v��]�<���O# ��3	o'\�@��,}Θ�A�!���q��t��\K6A-r���	��\�I ����H�$����aM���,v�����W���D(Z6��cu?@+�'���<t����c�[/2�rM|ǀq�W2�N���~L�uy�t�h�Ʉh�4|�"(���,� ��H�h!�_�y���@�n
O��;ęCB\���x��f����sE�ǋ��[G������
�S[@��t�8��T��V�H�������{|M�y���^}���p�.]�u` J�-�6s��~�*!���������.݉f)`,?P�|𭤜C�Թ� aON����Ǔ`����7m����
��G������gQmV��fT��.��n�/�U����ɇ�RC!�h���T��iy��Yk�aE��L���D�D$��H�/�^?c_=��TD�7�(e#���B�L(9k�S������w�c�{�<-���.	-9Z�jyn>2N��{+Fd���q��=U�}�oaʾ+�d{`8d�_�29�Sa�����<Q8VV��>����]������^7�Ƈ3��š~~u�ZN�	d��Kg��u �;+nЇ!A�J�H@nf�@d�Q�
4��������|pb�a)) �H1/~�\��eh�0��4�,a��}ҭl�X��<��/w� �u�әvVw���
���;��}�s�\�J�!`P}Ap�e+��K_�ؗG"sDކ.������J�mcl�0�_��l�m��������p�N-�����Oo��f�`�,%J���V&s���9y�+)��*u=3��-�Y;l�e�;(����q��Pt�`�j�ϫ��O�tg�>3v�֊e��I�.�sYT:��"eiU6���qX�Q�/ª������rTky��&'�j
S�QY1m���w9�R6��}��b���MY�@�S�39�ǚ .f6Ɠ%v濍�է՗�J��YD��L垷v|�G���3^r�b���c�%�h`v 6� 7�S\�ZV$�Nt����uq�7��ͨ�oQC��P���/J��ϴ���*l7���u @�VT����Q�� ��v>]�l6bց���K7�j�f5>M�d, �vR���'G�w�1�Wk;�t���!P>W� <36�Cj߃7�(�&���ݭ���}W���+s���o���h)���u�Ҷy���}���~M Hx/6��$6���c״B���6�@��.��꧳�-�_}�}S0e$�y���9@h� +���^�����䄪������l����W���`����]Q�,O���1*X�%^�r����L�{���]����"�ɒ(�mr�S��L��R�:�����-�w��ڔ��ד�Ü��T�w�F���c���5������j7�Eǧ���:�7]��v��S��d�>�h���Z3��P<��Xl�hH���-�$(�;�(�p���("�xCe��ݵm�`XS�?�ܨ�K�д^��2��E�<VB��(�1��͵�jm�_;@)R}��Z�E�3��rÑ�R���C�'�P����z%lU���5�ܿ��4�U�j�$G�����,4X���g�$4�N����F
��*c�*���Z��.��I������#A��4�6��g�W�;`��n<��n+hx�T(W�-�w�_�]ytV3k�]��rD�C>��ܲ��rv��ń�K�>�c_��G�$�?ֈ�6\Ar�K
�T������̅�h��,P�.*kj�r��%d���^�7 ��X����nA�5�%�����{	y8ɟ�u�zW�)>��ᢪ���Z�~��e�t��[~���K:Z���1�h3b�it�c��A,��4�9a!*V��4��ߗ��ӨC�d�㠡��
��MF<���B�+��i�G���9�yI�BY�:�������A �����E��9̥t���&��7~Lj�FR�ݿ7G��"�mh@A��,y��\���R��FzSy�9Bab�sR~+���7��tW�8�uI��8��8	P:��=W
>y�l$?L�������ε�"s0(�pWuң�1��2y���&И��8*p0ytl�*,�!�+. ��%���O?�-�� fK�Z҇_�������9�G)�$.�.�A��F|���6�x��5�e�>@��'���L\H�E}�,B�x��b?^����Zٵ������Fqo)��Y�����}����k��X9����7xrM��RE�;�~=0��ِ����<�j���H�q�>��y�2Hn�ܷ��]�r�سoa�`��[�����փ�nH�}^a�	��,���걵�쵻���~0�l<�25Ga���{�.�+��'tTb��3=n[%˷�iɼlQ��^�K���:<sv��]7��s�%�Q
W����-T��L�Px�&�|��M�]����h3��M��'��3���T��:H��M��CȔ���)>?�VOwg-�М83��hf�D��e_,�~��ʄWt/p�CJ�/����&��f�z�;�S����[�����5G`���m=�O�!�k���)1Ȁ��Z?�[��^�/+Ozg\ʹ��r
���Ҳ��v��.��&!_�]��+�a�6��i������M)Bt�\��Wȭ@�е2?R;T��ʉ��ɦ��_u�B�$L�Y��:ٰ�3$&[��G\Ga��B�S�G���3�D!�q���	&�Nٟ����Uq(�Ԙ\�!�Y��	�F=���H������x����Vzl���<��ə��+��|���@/{2>��X	�X%�J�������pE�> �A�{��"�}�������6#�#R���������wK��I���)�B���2�]|ř��F%R�"�7��tXyf�0h��t�j���� e�I,1�#ķ}����ÈL���d� ��W4e������)��ck��I}�Rf�&�H6#��]<-������1⑞&�cb�.�Z�a��0z�3>����Ӝz��@�]�>P�aR���XR"oMK:	q\��J�[�1�Յ��ȢwCհ@S�S, �>���8���]r/Ž�����2���e��X����zj�-Ll�s�O흈������
9*�.k����Ɠ��C@;D�;3�e�\�bĝ�a�&�vձ&�"�40Pf?�xT[';[����Ys����'P�7�jDy�U����X 51��"��O��up�xGDK4���ڒ��C�3@=)�P0�R�M���bS'K4��\�k�j��:^��VZ�	p��t�=�'��x��V�{���C�]�>ta��0I���Z����0�j����mŎ�m�p��K������{�M!��-�����Ji�g��w��v9t�����e{^��k�d���I�\۽��1��J����M��lK	-�O-��������m]fl�Už���8Cљ��e�_�/�d�z��ՎJM-Z�}A=��c|d������ c�}M`�����֎�<	'm�,�H��״W[�J���h�(m)M�L2���S�^g`���_��!6��o��nV�0��u�� �O�[���n(�M�ip6F���D
�#pw��֢�{�S��vX)�6���ْ�z+u���A����Ӟ�� �QzdՇ�D[��*�J����Ҥ�ǏI��а��tô�2͙�d�"� K��rZ��>S�IS[����W0�Ŏ���
9dI��	B�����y�L�	�O^���+��ڷ�������Ѵ͏�c��8�H�:�E��yq�8?�?�2#U�X��6V����b��Œ��� H$8G�+�h�I1A�1n'��+!e�뛀"� @ו"����^1�:>��[X���^	�T�.�M���.Ωm:;����f�HWG�DMU7F�9q袛�b�J%�,�!���#c�;\'��4yX���~/�+�z�$�ՕZ��2ri��C&��s�b���n5�/D�W��ˤ�,�7�چ��:K+ �O�N�?�|�-�B1B2�������']ca��My.n46�̌�3��q��B�َY3�]���J�"? `xt����[�	��{���is�nUw�먟�t
Zg�� ��_��B����9ׅ����ʟ�۲��3�/W��c��oz��z��� G�w�D��2�+�dKdׂ�_�=�5PB#}-��躌X�4�^��r���d+�h5�S/o$�&�,%�`D櫽U�C9��Q�g��8�EoyT� 7W3�-1���Ϡ��G��ݩ��j�����}���U�˴�!J2�M3�����H�K����2�g����gmދ/)㣄ٷ���	s��!ⲦIm��I!jܞ8�L4Y@��ӯv/�ﹱe�:��<��i�Ҽ�ctG Q�ttB�M�?�H��kvg�c��[h�:d�_c�T F���1y�"d��L:`*vՊT,���%#�rA@����o�e|�A�������](�P�/�A�β�G�J &`�&���^EuԲ%=�,�3��	b"2���Ȣ��ק��ф3;�)� �Vmݬ8c��/ΝM��Y|�!��y��%w��e�V��:��>��x*eL��(	�bm������͒a)A�T)���oq{o}l���TĴi�v\=S���ns/`��_����_��uͺ)�dlr����m~�������� �*A�4(A�_Jס�v���O�Ǒ��u��)�\r��}��QA1)���T?�%N��\S�X٬�4���gp�45!V����S�K�bo<|�S�}��˃m�8���&���w�}�kz���\�Cۿ���۱�PZ�gc<�� ��!d?��`��# M��oq,�x�>������+��BL�ڒ�Y��{q���q�\�OۮE���ǯG�}C�Ô��d�;�q�j]�!���&��)re�칄����{��֏��w8*MW�Q�d�K-�0�j�X�$Y8t^4H��EY4.����ʉR,�.A�1�<R��	�q~݁�/�	��B#���-:��Bzv�������q�φr+A����/�§W4$֛��Q�N
�;�iK���q��OZΙb�4�=��lB�B���ڇ�������L����݅������t ZMH�)�����5/U�k��Ϋ��}곹�0�5D��f�=�}� �i�}J�n�\J��-n>td�5�d���[5hu6����HZLL˦��mlT�:B��!�~{���jOa�o5Vc��dD�~dY��� �F�ږ�E*.���2x&\tG	�K���k�� 
�~��ϑ����fwg�`G�sLd�
�fFWz*�LU	�� ����<��ʿ䢔6���~C�9���C�J��zUi���w�|)���P���e#��M>�O2�L��\Dk\mъ�I6pT�j��=�>�����vc�8�=U����c;F;��������g?*�븠(콏O�eJ�zHi¦�6t\��AZQD:G�����Au;7,*t�Cw)�5\�H��R�ud{�c(~��ѿu���l��9ie&W�ϒqnV�Q���/~��]m2t��t'Wr�E�����M�~R`c�
�|x�	/15�He���#�� o��F�Τ��ssd�޾�`p�t�ᨎ߾>I�6�w%F�W�ն����)�'P):$߲5r�_R>�)��@XM�����Bî������wp_|6E2��ogi�����N�7�����2�
�NDvG��0�D�E������ؔ q�|����P���z�G�&Ҏ����:t'��7��3]hj�]��B̓"��V2��{�;p�|�������Q��t�D3�¤R��;�{�}缎�DT���'T��&(�l���ڇ��Cd����1Rw��k�����có!��>�=$}Ov{�϶�Q���b�6��"#c�|N��A�dk��nźHg�z_��R��O�e�'ve�N�Y��n����\BA����m�(:��fs�m��kgW� n���:R��'Ҡ�jK�G�#��HԬ��N�@r�-t��N���i�$��6+_��|CA���L#�����BNk�tҪلU��Y��w�]��J��k"�ܚ]�ߋO/���٨Qgڿlr���	�w��lQAސ���Vqؙ+��=E�����ߛl��h�Ø���p�rr�$A�L�#�PO]CS&��(�����a��޷( 6 ��2�+.�y�M= �P��Q��)��\p^�.d�Bڹ��:L%�{kh�_�^`-n|kk�(�\����#zw����gP�"�o~���� $* /0�u��J��x��_��^�<�To����A Rp�Jʊt4s��19 ?���Q��]%��L��J��c5N�r_�OQ8�Ѫ�VV�����!ػN�3�Nc�5i�V�)�4�cQ�p1'��̣��8(l�W�����F7,y����)��]�(bAڿ �3}�HG�~����6I��
