��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��?.5����
�(Nw���K���ۮCd+�>A)A�<�����i�'C��*����=F��-?����n�������T�P�E��(�z�)�Q��%y��%p��j�|��m+;�����.�˷��۠${Y涉��ل��5oyh������gοu�f#ව����E�L���a�S��L����>:ݳ��X��d���wm���6Wl=3�#����/Kj5��.�m��j�-���6�m�ǀ,���Ѻ[}�t���6H))�k" P,�_�y�l�T+A/�k@t�X�l�.��Vp.i�DY;��-�R
���MUM!~�g���l�U~�O��]Ҡ�TM���
�k?i
:�m�`M��$q�������%>�cҴ�+�����{�[֛��T|ս�)�ߑ��x�۲��U�����"�Û����̾J��ܜ:L8�+���|�3��B֍�5�G���&{�!��i�����½B��X�n7t�x����t;N��g���C�'�F��A$��a>��%���L4�	�.3L7��m��2nC�W��␪G���� c���$P�%���':��.iJyfGgOp���Xḧ���ɔ����i+l�m]'6����&��\�n�%a������,SvuZ��!h%���ѳO��=hL����³%����`&���&(��=4��WkCl��9���6�_��C0��1���6�;���Z�:C�"����~.��Tr��*�2�{��T1Դ��6�I�`����o��o:#�('�H#M��.j���%zX�s��3?3�����P���y�l�N�)3*Y���5�4 b~:t��
�3�"�!��*Ͱ�R�U�GT�\s�U3��<{�����@;F����"-�3�n���b�xk���+�l�����`ve���T����c.��/��l+XY��R�A_��`2}	E�]�]b6�_�#�h��J�gq�����9��XǠI�������(���0�f��>Ȗv���{��7��6n؁"�$�C�.%�e4ZG���5��~윐���Q��F@��LV��Z�~ܟ+3fD��E ҿ�IڢH[��1����ԧ�-8���'kϋ� k)?����o�d��>�s�H�a_�u���L����!�����<�.���;h$A�A�K���D�����tM6��	� J;0�����?��*��'�T�Z�P��w��=NA�$��7fIV�����&[T�K:C�+���� �![�c}�zz��������!3U��4i`v5L��?u.?/<k%)Zp1�.L��>!�����T�Mߣ��F�r��C˗��G{yA��@�E?�;[�$B$@&�����D�(]��j�/�	�`�~�H�ʶ�q`^^_��P���k�J���!\^�=?BlVJ�Ni����-�m.����}�u��J>��͝��5.F�����?�za%t�'+K�H.q�*����+�$K}��"]�iS���-`.�L�6\Ga7'B�vR$�q�ŋ-�/X�E�&4�1��j�W�b%�!�[�ҩ�:x�A�O�-|�`�
eh�>-�Y��tV}؅��I�{kO�H��N��Bqj�o�8�4BXC��7��]gb%Ն�	R!y[��_٤�i�-A8��UU uyA|^��������b�1`���B�@�8-U�\�H�d�1�p�@�w)p��zs�]�OxP��1L�,#�˦��e�������jk�豭��zlq7Kyׯ'qw>�D���˾�o�h��O�Ǌ�rб����~9�Hr$z����=3p��Y�0͸�;<+�+67[������ą�z�Ӱ��5�#D��z�#�iz��b2c�.>2���_͐A�C�T4���`7�J�#��u4�ӛm
��/���������ae5�1\P4^p��ռ��#<�q$�q�ȩ'��;i��Ц��Llv'sB���w�n�)�e5Vw�1�������1 �l7)A`n���$����z���wyZx�i�0�B�S���[%����V̫��}�(-��uM��jyo�؏�a"�#�ŋ2|�>��V�ը���>,��MN������8��4N�����=�\��HF������F�u���'�����*�^㒜�fF�T���ˀLJZ�?G��B��?<k��#iOE �g��b�.��` ����b�^8��2�����j���]6�h�����*D�kI�{̞�c�5S.���_B�l��N��v/�v��+����sױ�:\�*VzK� b�����w�7C`=�8�.M�ˎf��6s裆�[��@���V�3�홝Y2@�;���f>*+w����j#���ޅ<<S�5�1����w�������#o�H�����!��N$��Fl(��p	Z��w�.���v	u��Ɖ߻��S�b}ۏ���%���|������5�Z
ŠI�"\�Ҵ\��}� .��8n��]M��a�V���Z�j���J�j�ۣ)�N	��������3������Zn~?XAѨ;wI��9�t�Ż�&x�̚'�u�n�}z�\u��A��u�Z��pr'}lAӦ�#)-�k,ͤ:������<���|�(+a���[)Y!b}G˻Qtܚ�p�fzjò�w6]�S�"[�u`�Ӿ��
)�������O�!QSo��#[�΄�Zj�i���veGM�=�v2"iC���GB��}�n��r(��UR�v��Lr�&y\��>�X��E���ǒI��3H���'w~�	��a�-�>��F�*�#�] Y&(g�jpϪ��"�S;�ilJ�2�(z�o#-#��'j�ࠃ����!���Qח9 NI��y�i���wnQ��X`�[aS��vj;j%��r�\ƪ��) �"��$�Y��O9���*\H㢌]�AfJ�!���]�L��D����T�ͳLXp���O�`A\�)-�Ӻ�*ϟv1b�&���'�#z�3Sl��fA{,T��!X߯�Jf�y���g�AX����� ;싻����	crSz�^W��*IF�	��XN,S��QAa�$`���/D֞���b��)\plbRcLw�oY9�S#�ݡ��ީ�f�L�m��h���Y"o�t��{F�B2��Q	 Y�4�W����rDV����;�묶�[�5b��+��cԮ��&Og��"��*��.v֡lY�<N�`~XU�e_��@����@p�?"���L��߹�������j<_���K���6%`4+�\QLl*&���;�zb(֜l�E��{wfT�����xR��?���q����d��v�l<�N��%�sʆ��/^e!1o�X�INe�*���(6Yo'wy�g�k���7x�E�<�c�V�KW��g �(n4���~+z�ħtam��l�T2i�!�*��ca�8�f��,C����Jx��D�i<�?M 1���z��\*ZP}�w��`��賖57H2�3R�����v�[�mt���؉1d�|6� %v���H*���>��M�Z0��	ţ����摳bÎ���6��<���^mn)�W�i��E�А�/=j�w$v���
*Z��,i�?�q�k,e�ۻ*65��¹�V�6��Y�֔[�}XW�#�O7�t%�%cwE��#Q�Ln3�p�*�<�8�`^2I|��W���Y�'��/<�/!Ǡr�_'>e�A�����wG�P5��"f�M�Y(�鰏��O�X��@Գ�|BP�C�㠙`/�(
��e�oH��%��TEA�t���n@Wiw��_�x��0�-��!=}�y��3>a&ѓq:��c�0o�B�#`'��n0k{
���|�7ϙg�s�]� ۰��p��\I���=��9�W-���f����Kv��2���?:��[>�y�`�;��C�F��V�#CQ=�3!���4 � ��Ҿ	��Tں�"g
7L����ܛ��Tq�m5A�	!�ee$641K���E�����P��dER��dV��{���(��1*ˑ'�>��@ �Q�4��&Q�N_v��!Ztl��s2YS��֒��p\�ZX�6�u��/�/�S�o
�ƀ��P�3V�U��C�I��/u({4�p6XY��k�vn�y5��(�x��ih�����\eJ�n<�����1���e1�]a�J`zt�R����뭁\�a��Z� ' �/O��7֌�D��ѱ_l��n�m�;�E�$�{�����-��ɱ�S�a�Ů �j�F~��ӫ��ѽ�n���+��۞�[r�A��q!'y:����M}�]��w���U�rWmv�A,����N|����sVJ���'��X�)Ɣ)���y�Hl1�	�m�V�D�T�� qe���m�t��g��Cd��%��oQy7^+hz��e��|~�@�7*�:����� }��_S�g��yqxLJ_����P$T �iB�۹���[���b��H�9��瘲K}٦�A��a��9��e�^U��{>L��Xd��o"��>����0m�ŗFa�n�`�wQ���rR �J	�"oY��J$>��e�N����g|��1n��]I��ʱvj?��3�)�37w&n������H���۠�C�7JK�����ɶ��A�Hm?[C��#!��Q�G�T��o��y�d^��и̰FӀ�hC֝�|%?�Y:����S�5LC	���xm:�v���B��D���v{xTP��U3ܦ9�T��Ġ���/�g܉g���h�~9��oy�_�{c��8c����2$Ѣ��oR{���v�2�7�a�I(P,��#i�z��������.�?�r�/8�X�:`~$:�k@�0�;���H_[�J�EU�Qr�n���}�j� �D��1�p��$0|�Jo��X�w���n��td�6���I��5�{���_B�,Gc��������۩�n������b_����E_�b\I��l���i��_�C�zm�m����FZmu �m�^�"�z%ǈ2��~a�o�(X'��E5�0OԾi�'N�7�2��z؂������(����%A��td#�x��g}�95H�>~���C���l�������$q��02v��@a��7�ϥi���<k�N�����10 9�s�ˠ�٭�)�c���@W'
U�5�+P[�w��*7������]\g����8Ll`�H�S1�5ò��DZ&ƞ�5�R�p_ �&U��Z\]\OK��5��_찥
U�w�4�]�L�����" ������j����dl�3?��BE�5��ӟ*	 �g�a�CM�&����,�U8��9 U�ORo���+�@�"	�Eu0��$�v-4˧�V��x�P�.�X�u#ady���q�|�-)1m��ZcǇ+� �Fg��F�A������xɕ����|Q���7�gc�n���:g`9B}Z���QY��C�a�x�xb���8��gF��̖{�m�M�K��~��nJ�QڥY,��6�y�[:��ڸ�@F���W4�89��.�EK�n����B�}��V�X��Ez��"�����ҹ`c��:�H�����귾-�Er~��b[���z뀰��_�`$2w�0x��L��zM��2(N�7oy%n�����\�ۙ�z�����h�>Ƙp
6�B�#*����9^TL<���O)��0!�]�,:��I�l�/ֈb�+^H��O]ː��ɳ����:�Ɋ�	�v�z`���+L�+1a{|�壡�
+9�}���dl�w��ﴦ}�
��
�����H��׼���AN=�Goo���\�S��5EX�W�a�r���H"�Tz"{���9�t<Z^G\Fu��
��s�ǭ��3T��"Ҿ�e�g��F�_�͊X��#��X�	1�_ �f�H�g�P��;�Fd;}�T�瑈�� �e��2�ڌ�����s���Pg�N��w@��(�&����g�$�V����ʟI�B,v�q�D�흑f��ԋ�W�Q�������A�S߻������:�ƍ�y����p<��L؞��vm��������8������H*<։Q"2��a��\�*�7�����2 ݞɤ�a���2��㢟=��)ĩ��-���N�fwfc`�R�9>p�g�T�rg���b���:�C@{�u��a���=����.K���V�ȕ�^�kPe���<��"�M_��L�M�.�(�`��.��h���Xܤ?��	�W�mw �0Q�;aΐ�>��\P6'��oKh�<]`�NBQ��̉�>�p��uQ�73�8'A�����er��X�+�6�c�~p	�����Ńe��������(��c����-w�ÐaS�Z F�}��ӚGs	��E�vVnf]lP�r�s"MQ�>�,	zy4�o0R��G����R����
�Kg؝ۙ��V�`��|���|Wmd�X��T@�? K��p��a�]p����<��{�,��5Y𧃇k��x�;/�\�ۍ�@�
�A�Z��Ɂ�2��� *��Y����S�R������R�m8/���^��kq�X�[	0�VD���!G�{�2���ۼ��}@�gPg���
n��A!�g�Q\��6`��pu��� �g��(Sf�� ���Ӱ��l®+��
�rI�8߹x'�}i�QZu�)���͉S8�-���xnفK���Ph�Y�L95]��/w�h?]���\���-$�-���Ħ��L�FQ�M��D��!�12,X\���Z�m�l�ĆM�U�I^v
�p~Eb�T������-S[;��H��v�ˮ�u���9<}"=�GX	�ZZM� ��`|]����x��=盿q��q��J=N&⠊��ר.����7=P��ݢb���<'>�� �I��	�lџ3V�,+'B�s~��K�������D2W���U<-�1����v�W��BS�L:�Kj�,t��4�NB�d����i	ˇƸ�:xI�:��_rv$&Ii��	�l���'<o��R�>酴��ANM�=��~F��eCxP����*mv,�J�]{%ȕK�f,ů���NS�I�ykjT�nt�����l�7`ɩ[2�e���dL�2�::D#W��Y��t�7�'��������0˭8�0��bi�(}k�Բ���d�+�2.�{_�7�e9¥��A�rrg���3x��X@�S-ܖ�}%��1�����~d/����X�U����H�I4�kQ����+,�z
^=Ǩ�?�<3.���]���tQ4�;������[N���޽t*]o�زH��j5���g�ݙXp"?kJIxZրP�hV&� "�I7L���x��ڄ����z�R���5�Ȟ'y�+��X.��(��Cy8#c���w�Tp2��t�s�1�a�'Q��i�,몜Ry���럦E*I�w�2p�����!X��|^D�n��g8ń��.���pm��t"�Dgo7�U�A�h8��Ũ&���k3���m���P]z_�nֵ�{pb������?��T+���;{8ɞǿ�|.�7�zo���Z�k�`�wCo��I]>��o4h�c<�NǣE�Wݷg����|��f����.�^����Ck��V;����2���[��y�w�<�O�>�����hy����9�8n�>vm_��Z�Aȶn&�g�:ܪ���T)�ы�c���X�"�lN�0���iV�J5=J^�hAO��M�G���U��U�^G&��� �!�a=,0�u�d���ۯ0j?�.��<���AG��y��rI�ҤX�^aVqa���1�j�5ϟ�֚��F�Y������|no�� [�Ʃ|ݧ�ZHoo�/҈n�w�1 ���۸�!�~rC�����om�ˢJV|Skl>�?xig�U�Db�5��&������ _U��)r	<��풹7;
 S�B��o/�_=$�@6l��c�>屢��b�7�=���'YS�����QHJ�����&���5c0�Ë"&�̋tK@5�&��@�!���Atrem�å#?"_k�w�~�����K��M<5��Z!eϼ����"�Z�'X�{o���֙.V#n�U_4�?3�٤p@U�ױY�w��g�5��\D�Aɵ��4��ؓ��W��@����ؚ� ����y0���i��a�A�n�H�+�8l����p�ˀ'���&۹E���̛Q���6C?7a���BK֌�İhZ@�)�a34��i��"*����A�i`Hj8Mp�d�۟�;�n����V�S!�j��/Oqz�u��QxF3�xVA���o!�Z�R��ɴ��S���!$R�s�oC; 4Yo_�����d�Z��Aߛ�"Ky	+�I��AU}�`��\{O��k�.�~�ќP�̱�:�zػ���)6��J�khE6��rQ����*G6�����0�ZV�վX�D9?�~n�N�N���f��ĜZU��n=�H���"��r̼E�8��vYXl2�n
n3����ئ��(Hn�`M+��*�i��( Ә焂;��!�0����S���	���\��:�V罠���օ���L�fN�sk��,�V9��"�E?t<gX<G#0���7���!(����������w����@���t�g�������$~\U�.׬�����a �9Ҧq�W�_����Rh7*e��߬�e|�����Z����G�0VFw%FH@���հP�qx�J�����p�#q���T;ǃ���I���{a�Z2��ڀL%�C���_#M���o�dS��c%��USd\C�wZ�I��
2i�g�Gs���J�v��Ji��px0���~���\���@;ŕВ��M����q��|E��F/�n�\P�LH��x�����L�McX�Vo	�����P���o	}�j8@$�`����&�P�X�� ��2V�m������3߸o���}����ƀ/���J�ʨ�C���]x��~4)t�T]�>�,H �)��N�DV�y��{㊯܀̳����#jh��~9+��A��4~{�.o=l�Mu٥u	���RI�ՏUI5����`i�r�&+Y�T'⦦bY��S��0?d���*��$l�r1+��S���,����G��	�3���NJ�f����rzo�-9��.��:_�:B����0NS�X0o��:6�VH���C�a�� ����#GG���U���֐b5��RRy��\�ݣ�*�x4+��ݲ>f�GT���"��V�]y}fe�<Nfkܼ�t�2��#��^�F�������U�P6a�d��o�sDl�|�xW���i�l�HZNA�Ս����Z�-�z�C�d� ��bx[���<�ҽ����Σ�4�yo%>B�[�z;�ոY�>��s�wᙫw���/Y�d�t��d�:�Ϣ�h�����ч����ߝq�v��&b�ci(<��`<a���jqH�]�GP\	�y=&h+�L ��R�QF1RF���*�`٘oG�0�-�d��^D�ܶ�%%�Y(��"���B�쩋�8A��j��ݻv]
Z� �t�F���Q*��0���Z�P}x���\�AN9��Ia
(a@�����\�kbc��Ͼ��3H��&\���O�#�Sp��4#{/i��/	,�(a�0eY����n������	���/&i�l��\�V[-`�X�cQh��?7��r�ZU���)���cO�y��)B�4EkS�C��/<�%���ţEa'�r���L�w'�g��Rk%�����E�����}lC�?��O����v���1%\�4}�-�o�t� +-�7��gJTއ��g�F3D�M������`	�O� ډ�����K����s��Z��� G���l0�E�A�@�*�'$���X��L�՛�<o�^�,� �k��R[��W�r��&���@�nk��Wm��y�3D*C5_Q�ɡN6��}VQ�����_�V�BWZo����t��ï����c����js�g���6դC�g�ZY�&|�ʈR
D��[XD<u���<llb�Y��}�6�0�ӏ��e.���2�j��}G�cR�o���{������G<�&Z�(Q���6�O�L�ֽ�X�HOP:�dI��\�P��{BP8oG����M
e�P���
,�5X��K\zP"��F�O���০��M[m��@��6�BF�Պb�=XcC��G�B[��nٷ�FT��|��
�1��g�C���+��_�C��9�1��>�m�xzI���TR�� C�+�5�`R?F�F��Q�Ǫ�O���9������H��=�T"'�@�v��P£�Ic�Y'؁	����ǌ(57]+O�?���sA5��,���^~��X`�X��$�8�:���8���I�D�[�>%�<��\c����Ɉ}�iѻ�f������| ��لŋ��H�(dg�w*��=�р�y���@n9�'m~�ᮿ`�U�ap�*0�̧0���W��m}�\Ac1��~���$�L�����	���j����rY֬B��I��7��Q9�H0r�K��[�H���1:�W��a3��nИDd��`(����!��Yǩ:#ڏ3"s�!��uy|�`����ѱ2���y�9�&������A�N�	L@M�X7��q��,�v,��e�S�yi�n%G���g.-Y��}��?�33	��=�V=W�I�ph=�����|�����9�ņ\E	���0̫:ײD{����DNUSwa�dk��1��%z<%_M¾`�y��8u��tz�~a���H
��+K�L�J)�����y5�rNԊ���`8��8�
10>$�z�5�C�<������g�ޑ���g��П�m�쌛���
�!�Ȝ�I�h��b
���hy�^��*φK�����������+x!�[%����Y}�='���̀��&���d��5�=��eY፱�\��9�Ī�8��[t�Q�:�Z��]k�����ky���!u�<V\�!�|��~{,�Hy�����/���J;`��J�n�+ U������n�oa0���0ʈ,
Q&CK�~��a�68/�)Ȳ��)l��ܬ�Y�it��}�ڽK�)ތ�mrr��/�%',W�Q��/˿��:C����
cTM%�OA��GBB70��:!#�X&Ֆ��v݇�Rm��G�9����}3�)��hJ���ޙ~}}0[/��E\�)a;>w�����@qI�~J�}}.�@��]�=#���C"�_׳W��w��ҍA��s���~Jv�Fj����[2��t�����<�F�<B�oкڃ	�2�Io��9q2[��Zw0�a' ���$M7dY=���jB@�r�ݍ�~�`SЧ]��?��P7�������;`-��_���6)�%��l�U^KCV���	���K��F^��#�O�X�{�9}9�u����P �������4yqX��p�B��T��tM�jn����Y{v t��3mH^.��Ʒ�^�HZ�C�+�_s��QмD�3�F���#�_t=���6Δ�����������V�p��Lr=�ːl�����4��̧��3���"�_hӘ�q��%R�|0��B!��1���������K�7YK�+Х���Z���i�<�Fs���YE���"�� 8vQl����-i��#�����b��D0�i�M�2z�Șӵ����>
~��~�J:��ه	>�ޗ��.$Eq�W�T޵H���>F�>k����]�vy)(�w���I!ݍ�CY'��DFu�����po��l���0�C��V^��Q������w3+212t�4+W�{��4˶R�V5p�O��Ϯ%����*���pQ	��s�! m �zR���)�M4h��V���]L'�� CZ]SRC<y�v9������Yz'�1�?�=e�k�w^;�q��*��]��������G�m�3v�z�4M`�?	;j�B���v��;7�-�܃�ȶ�
mZ|�8����)�Q�q�io�g� �	�iV�+��z>�>�Ӄ��c~m�4J�X���s���{�#>J����-��e
Fj[��_i�����d?Bn�d(���1\^i2,!���qCt��Jc��Y�M�,�_lτ)Q��e��4v�������ۀw�?9�/F\����<��0iZQOq(�ѯ�^�����q@EJSŝ��4�$z�h�!4²�ֻGFh�0}�=����'�y�����p�e����u�ό���U*Hm��vy�9�HSս�춉�%
o��x�IP�C�x���=�e6n���YIs؝�jD>�2k���� ��('R����T¢������t���:��X�����Q����`���� �6����	3�$�w�M�&���9�[�JN����.��`�]B�C2y�4Xj�3���+8DwA�2|w}�zrT�B*�%�e�	KS �
wX6���+�M�[c~��qV��b�
\��;���eb��C����m��@b7@`up��-��gM�Xޚ=F1�U$��Z܎a�#am��f��OY�]�1g z�^�YУ���R�v�������!���̸�k ~�z-*#�O��
�I�@�s�y��t�H��j���`��ib�21E~�����A�i
ɴ1�D�u�:�tŢ�H���.`|��!�w�P�[��������m��y�;�g�ǡ��҇���I
R��E~����Ȉ;�|�*����'����D�K�^~���^D�mB6)�JؓB?�>#)NO�I���,�i87��9�"�]�+��
�A���cY7�au�	�k��Y����X���!L�+�b��-i'�vNn, ��2��a��K����ȥ�YXk �5�f�ZtoNP��Wtţ�p���Ҁp��Pr9�6��\��)3��Y�3��9�)z���e{��޴�ꄔ'�jp/�4�A%D'��ı�Hߩp��sĻj��/J��Qm���R|z�UnP�|�/�0N�A������PE��6���ݪ��$t�B�����W�n�l�N�N�H�'�R��-w�����f�}��?%�A���	�=\�K4��yIznO��łH�����~��O�GicJ�-�z8����*����3�ڶ��׶�'yA�AGZ#�h���o
3�Tx����E�L���2:b�(B�5��7��7�2��������	~q���D��'�{���"��~�����5�T[�� �qj���%
���hl
`sטG�@nDK���H�)��Eu6��y���S|��;���o�ϸ��؞A�F^�9��K����g"���������g �����@TqE�1Cr̩�(�Cۥ���A_y9�Z�Ѥ��X�`59��gA¬��|������=��	S�S�t�U��T�Y�sr�&I�B�ܴ��e걢�]��6�ύDi9r�����Df@��'(v�]�q��J�����\-���K�ы8�0��df�J�x����މ��>�>*������1`D�!��/x6��gr�m���P��[��L�v
Z[���a��XT����S����m�i�J_�NL���a$^�wC�a�vc�|�`6�Qg���,�q�2�Ih���[n��`�QG��ԇ�&��"��|0ROk�-�r�/:{�O��B zAs�,��'3�e�]��k�A��v~�Ќ�0���w\طR�	��b���+�D���M�Jwɧ����&M+��j�Dt�\W�h�uo[5K���j���W�s �c�i��Vփ��-��'3��xj��ں�N^���*kl�X���6���QuK��᪁>D��ю�����}	q�{�߅��a��Tb�,M�&
�p�n���<����֦����Ƨ��d�!ߒb]Ӆ��J��f����0�D���4:UN�����o�~�氶�?�?�Pl`h�B����g�͵i�!i�?�A��I�R��'�G*;����ꏯh$�"O� JcU����K��M����ִ����5FPw!�fS<���옏�D۾���&��ڊ�d��v;�CK�!._��@C��t;���]�k�� ��;X��MZ!��d�Wym�JqЃ�0y��X�~$Rnt���}7���'������Z�s!�e�Lcs��;�*I�>���a#��J���pK��=q����SVn�P��;7��`p���])�͑SdՁ��+���+H���{5?���pǘQ�^H���ی�,�-Y���+�z�Q������1r�ww��
��2C�������-_�~��#6>��}ǝ,& i�
�6C���G�1@�?x����]��t�?u�b�{�����'��w~&c��H�&7�a}d�F�~aWh��U�[9]���)1WD��f��2�
�` a��`/Φ&������@B��ow��B��T��B�O���q/�p7�¾}��{��i�<��}�\��PO�L���=$x��Y��6�+&��)��K�I<b�	�D�RyV�Y��>+�����J%�dxW�ￄCT�L�r���U�B�%�5�WO��y��,�p�9/�/W����Z�"��Ωj7u�'P���F���Ìc$yq��B��̭|�Om&�1�p@���.�t��g��RLY2�+�Xȑ{|;�zמ�Gk�8�;Ad�hqS,$�R����8^%�Ls�`o��9w}ϐ�d
���2�d(9��Z��W9�_S+��:���C���-�����-�7K�T���L����W��wO�BR����w��w������V�:r}��nO�����:�B�5Z����X����)0kz�V���g��v*�u����]�(6-֟�81�l�_��:\��E�N�Ym�-4�
�fKș��t�d��Y�u�}��7�����n#cʏ����W]k��q~��+�v��ٜ`�a�`�n��{W�A����/\�u#��d5 �=u�Z1���^D��ᆘ_]��̵/��Zɹ�����Mq����[c}�qҬH0�W`3��:�8�zϴkN��k�<���I���`
u�O�u��gP�ۓhk���eJ���H�L���^uעs�2�(�A'��x��P�����>�����l�m*�4H�`8 @[Vwc�.h���� �6��ߖ���ƥI$�8�!su�#Y�����K��rK'��!�H���z����������+'ex�0#��n�j�g1q�&����X6�LT�ۦ<��ūW�b�}�[������7.���BQt���E���O@-��Q��Sy�V��b@�ܱ�!�q~
P@m��$��L��EB���q�>��!v�AP���QC�����M�lbb2N�>�8Ey�>Na���3�oQ���$*� 2�ֹDwФ��eC�Рj�{�IO%��).��O��|�50��l��@�c���D�:LMύ��9xe��6�N��8dAJS��u�Cy�-��t7?!mRC�"fF���,*��e#�����!�<Ά(I?9Eu�"��ڵ`��_v�!�������rMR&O�� �532��ry����*��f�˸�(���\�K�O�9�����f�'10�]��5^��|��jS��:�J��B Z)r��r��Ҧ� 9�j\��5���U�K豋X��&7C��SPM�:-�f��'��5�Mf9:^'g��-�2OfG:jC����~MjG�^Đ�,W�W6�D�.��q���L7�,r���ծS���6�:��7L������o<U)W*L���F�	,8P{��Zi��ٌ���i���K~|_�׭L�6|@TX(��,%�h�!�V��?X�2�4(���]��]��C� �D.p�S�#�������@c��"vjc���g���B�`���ƙfVr�~�h�Z�h��H�Y�<�z�; ������Bd�T����ѡi�dY���Eusz;x*><��t��#EA�����V��l��-��"k�J���F��5v���w,�����_�(�MR����.o��bx�L0��CCҨ��J��uM�9����Kچ� �X� �A3LH�a��
Ƙ�v�(�20�x�����	�Zy<㵬��j�! �U RԨײ��p?���R����OA� ^������=q[�#}8X����d�5^&��|�i�e��Ϟ�,0�O;�c���ŗם�未?ܺh��O�}��������6f�Ç!�����)��C�u4��e"�S� -�⺜ҁ�n'���z���.���?@]�dfRP(~��O���(r۫�2B���o�1�����
-���UR�'Pr��܆�舣]�H������Ѭ�2Zz[�b���g���z����F�[kC1�5m�ikY���0	>�YݔQg��81+�F+Kr!sS!�\�������>�Q��!W0(����_���w_���� �Cȿm����d�O�+��_�q�'|�,�~N��:�X?�'��hbh���Q���5<���!�ǭ�������2�$?^�G�:֗�G��}��R0yi(jrIL_at�*��#1f,���>n|!���c��]X@����W̒�>?ם�e��q	�z]n�p�vW
���fR�&~b(b�:�.~����MEf���#d<7(��N�l:t�t2�)�Sm�� ˹���io�����S�$5S�4!��Y�؂!�0��GdO�XB��c�Fz�~��"�Փ5�r�E�/��R��X��$y|D���:�9���-�&�]?��
��H��/O�4���l,s��>�jx�D��U���A\mkf��T�ʔ
a���k�.�8�&�5f�i?s0M�V�"IgA�Y�y#Ɓ��x�c`�]�t�]O���{{p~�)�!:l@�t�|�w�i0���DV�a��S�:I�H��X������a�d;;ձW�.����n❃g��b����j��{���t�2p��6g�U2����_ 	��0#�d$�^%'y�D�N�|iX�4���9&�KK|uۧ�H��&M�P2
D���	SRsӑ4�dm5�U��me���ճ���[�˷�as^��͓vW��5FA\2ؘ�����6l�xi��!��T�� E�k,`������!��&�^#;UV��)1�юDc�g:�Q���W����p��mn��G��9�x
�8Xތ��<k2E3�#ތu�%�~?� �B�����Y�<���5��D!f���b�rI!�pj�C�z�Q/ ��m�a��b�� �\�FV6:���q�9��<�
Y��k�qŲu*߸SN��	|l�M[�i}�l�;��/�}��^d!P�-�)=f$@��LF�.s%�qNg6��l]� ��zC'���k�0�)4b��JFT���N��g������Y,�����2&�q������W2�N����Ez���ֵ|�NsX�>.�GC
7ڠO۩OQ�Yƍ\A�!��E�R���/�S"[K"��LI�j<�ᗄ�ٜ��
r����w��a�!\��$�O�q�4���m��-;�[\�'sڴ�?�MBb{� uZ��uM��]Y��!��7�Twe�o�\���-D[^�.cj�~���nhii?��k�כ쵐A��1����~Gě�Q��������0x2�|����C-�?����	�=O6���'�;4�� ��8k��& <3)�Dn��|�����1:ۗ���y(#�$#޷=q:>  ����ɥ�\�fzm�}��Q5�u��:x�.�Dc& v�ﲦ�)�kU��~%��~�����7�U�{�K�ڰ��������]5��aߧ�^@���i��`Qnl�7���ڂ��j_�u��8�J�b���(�/w8}m��ʆ0�l.b�t̨�:C�5��--Zz� ��=a����	�׵�O�T�G�E7V���ygX����~��;v���]�<�)��*4�1��@�gw��w���i0���4T�������>9ҰF���#�Bՙ4o�f� J"��MAf)�M<�g�J����v^��<�p�M�J������3�����,!�W�[�X��$�H�s��N9�|�KÍ&��l̽!�_�
$�q�)���)z��k�/�V���h,pqK	�%��������kǖ�^u0�f�hGؿ�w�@m�}.AH���I�����3���y��ϻ�F8�܅��d
I05�>���E���r��i/�������o�r�>��1TaG����t�� ��j�,�8R ��?OC�4��
��a� T���XZ_�x3����Z�WF\mw]��E�D��֧i��Z[������I��x:ʝ�f �gpcyn�)2�Ne�R莬pY�F�
�x���D�UN�϶�ï�����=��{�I�{\�d����C���� ��S�8u�ӆ��!��O�`;���7� �f���R�"�R�U��_W�=Ա�P��_h�!��ɨc/��8��>Jz�	�ov���1Q�0�eɊ׳>ޣ�*�z���6&��	�x>0��B��<��%<��I��&(���T��8G��`Eh��i��o��A�3׸<o�u��'b'h��"0�"�(9�	�5n�aBA�i����"�����A~Թ�.�\�`SA�蓊T��FK"q�I��S�M�i24#�� �$�-��(���L�w���[��V�h��
�~FJ�s���S&��E��YK�@+��`gκ]O��%`�`�ǖU/�<�-J���q�ê�*��?tN}3x?��q�S"�1� X<�f�
�b�8SODKj2���c����
���TN�ei8����Ku`�6�m�znZ
�hVY�n���q����7��2*=}Z�t�s/C?��GۖK����s�zK��3M�p����2��;:�1�g�Rk��.�C₴>�X�ܞ7��}`1��E���F�����5�Lq����LhQ��#�ށ-��6)��Iƅ�H�z����e	��H��*�����s8�T�y���4���Ghz@�#,�l�>N���:Z-��º9x�H�^�tB�D�3�#*&?�di>�8�9J?�_�C���D�|a�[/c��^V�/�����f;�찃��٢�%��|�{���y�~q��2����@`� z����m*�n����kj+�@%��@\49Ǭ��i(H���NLsr�I�Uk�*��H�t�!zBg��^!��Xȩ�=��ur�}� 6�(F�LJ��P�t<{k�l�,�	1Rk�.���M7�D�4���~�z���`��ш�w2��&Cb��bק}.�B�h*=M��܏���'�/�p3�2���dо�ǋ�$ߌ:��|����5���AX�Y~�Q�O/a>@K+���t�}�'!Z�ϫ�>}X�K��4���� b�����d��x�����|�N�j�x�6�������,���2���IQ|����bx*q�'��!�1�u�L�$��f�!�A���� ���r��gP>ɌE8[kk� �I�e,��ןzW}uF�j�[������1�� C^'(�Dc�UGZAs�ǣ ɯo�E< �d���lo��y`A���,F�p�텖߽ �A�o�ӎ<JC5W�SA�N~g.�����[ 8����V��Q��%��zǹH��\�L��������PGm�V�b�XPJ��b�ĸ#��B�Qt���,qҔN	$�&0ǵ��]�8u@�P�H��W/�x��i�o0�{�&
�lE�N��qn�o:;�E�3�G���ל�"�q�o�ةv����zw��A��l�(��A�������ӓ�D*�gG���5����Z�g�14��u*^{�i�ʱ�(̴�=���)L���4�Z�U��|�9vJ� ~ �x/�5��o����
�X�3�<��_�Y�~�1���(�s+:��<���:@�k2��W`*���:	�ߪ9���z��lhd��y���f[��)\�o8�(�lOsd�Zw��R���`���3�Z��?إ�����cH��s���
Ѿ��=[�ͲCV\��ǈ7��ͤ���?�+� �$�W����ݸ�@ǧ��y�N��:���Ġ^<����p�z�ۧ�{���xn�l�(�e��V�1�����?���9�B����-	���,�50�C\7��<�3���Q��.'�{�D���K={}�C��jO�۶	�b5{��c1�0��#V�R랽n��nj�B]�`QC���G`-�;������J����PK~��v�V���O��1�\w\ ����z$��r&~�5?�����q�͊:�C���]��.�a�c�O4I�7E@�>�5s�ح5����xmٕ�ɩG*��ϻ�.�&n��d���럇#.���>�"HU%w#GZj�$���D{�hq�6��7��>�k��ݭW���1��7�x�0���[�YD��ۯ{����ۇ�(�#P�p|,�*��)9(�F�RP<^���b�U?�ܧjH�Ӑ�j18:/�+�&u�>N6�o���.S�S*j´�'��J0m�\�i=ԅ��q�GӬ���\,����\�U2֓M�4��R�E=C�%>Gcn|��W���=nn}���*�u��M��O�;�Ƥ@�x_{��i��� §;�U&j��>�n߫��C�'k>0��������$F���I}�ّy�5t|�L���X�`��0��lȹv]�K)�� �l�����	<�K�UYS*��%8@��� "�.]�=�"::���������4k&zn�î����H𧓭��d^~!���ĎO���`u��i��+��P�y�ki����y�W:b���f���1� kv2Q���x����u	��r��ʥd��VdK8N2�=�}�":pʁ�d����J@Y[d�N�sC�˷�n"�����EZ��S�k�{�yO̰X]�<U��f�BB�0龷E��,����6�0f����7�3���7G���*a�ŊӖIL���&��\�kM�Ǥ���~���
��e[��!Qz/�G��{�WU�}��oz�$�m5y��:���:sK�	?�_���˘O,����3�)�?u������ 	�^�Ai����Z �Ӥ_���ʭ�Bj�D�w��
`&�ߓ	n���d��C��P+����I���-Eh���k���6�r��O�f�a0l���;�|�D(�xv_Q�0�}f5~���nZIH]C�Ni�]G�8[�^^�ݻ���Pg�Kq��O�q=���Ų������������E��y?᳨����Է��ێP��j		<dp���\E��dF����?;:��#�c1��g���� �����6	�+�ƈ\0_��W��-�`s�([�i�@D�]j��&T�֪�^���+���T{���;37k�y�c�I��>	5q�Ex�����?f�_s�����m���K0��k#?*�[�I#�(�[2u��i/w5C]-��;���]~b��gC'l&S�/��V�u�a��<����Y���a��k�/�i����$�Vm�q�X�9���^e��0K�N�o�Y�m��t�j�����[m;r�y�z-Q.::0"�CDƨ���(�)�v��M��:��6G$��u�A��B�	�]��(�42��K�_��nx�ڕ[G����#�1�p�Wl�n �K �w�y�f�Jr5dЃ�f?C�[ڳ��G��o��^L����[��Zr\i��Ո�/v!G��c��bE�{�ƍ�C�n�C4(�Փ�ZC�!����e��I/���K��ZO���A	laDMd�$� �k�.��f~��E�l�3M;Yz^�B�^�'��r��Mio�p0o���="��Q��l�N-*�I�3RQC��L��I
�ϵ�͑2#dz��/+�WlB}
��(NO��ry�T�ޝ=��|m�-:V[c�J�u�����La1��5��{V�iX؇���k��6j�5*��|'Er�'�g���|�[������jPR����ꈷ����i荀5`��)�X��բy|od�h�x��wIam�P������PbÉ�S����3���5�j4�� ���|����{`R�")%tm��ӈ!�{V<gߖ�6������,�YG�$q�5'�SN,���1����9F\�nx��9�S�~��������C��Iwd�^���BST���2G���q-� Ѯ�K�9��e��'���]�@�����O�j�@�I�xf�\�>�)��C�~-��ʍ4��)sfJ�F�a���T���!\Yk5Q�a���=y� �i�n����˳�"L]_y �š����A�r�+\&�[F��2�>v��Z�N������x��a/B�����c1|w�hč�1�o{eN��z!�Τ*o;=��n`Q�S	�����?f��r��v�M�r����O�+��4&��q�=�м�nчd�2�d��l�����<����<s����/0-	��m�#(�Z�%�O�?�F���4t�F�,�!I��8�(�57��--��SQ�`���~�yr�ʿ�Ij��/�xaE�C�&�3�ܩ��ﳮ��ݿm
����k_s[�G��ܾ�����Dk��n�K'�d��d\ ���PP�o �:&��Sڭ�Iݣ	c1����y���o��NX�!H<�)��3d�琢�nj��*�b�`R5�����t���R�����y����緜C��8!��!x�X�yP�Z���2�WKqw�C���Fc~���<]W���g�IFEشȃ�װ���2���cUi��b�
��ھD�E�l�1įOlL��K"�sʓc]{��F͵;��y9��(���v<
�;8�Q٘9DU�3U3� P�À0R���XIǫ�J�KC��L��/��wz@e�f�*/�I��4��6<A:��Z�&�5�~d�=�2���O͚�����>p#ζֳ�� v۟�̰,h���A\�\�r��h@d��T	�m�;��5a���UmԽ$
��f���*/w�����W��i9��3nK~Yf��ZuNC����t�Ir&��ƣ�)G��] �\q�@�|Jߎ���0D~r�FT�pVl���5A�^2YH�⩏�~��5С��U����.�����Xۦ� /i�0#������%�y<�0�C�l��:{v�:��j��r��[Bu���J�>�@�GIȁLM�<�ocF�11��e'�q법B��nw�z~5��-� 9G������B�V��@�8�$y�r
�>�e�fg�v*�j�£���-z�P�9^	��b� ��0i����u��)`8g��R�p&��u�����?z���@zŝ�l^������*�z�3���}�Cρr�������KҠ	ڇ�M �aǀfF�IY�Wt5k�B�,w˱����T�
l<#;�������	L�d�`N�������!sA��\�@��$�wV�Hr  ���%��Nͩ�Ъ������-;���"�xx�ś�_�|�=6�w�
�O�G��9��J�|t����@��R���*�&���+�C�,�F�Yf����� 0u`��[�Ȧv���f�^G��l4T*_gL�#�!���"�X��V�N۴Q�T�Lw����H�0K6�M��F(%Š�r���^`��4���v-��j6�ȕ�m�� <�8p~�;�f�G(��Е�4AS��5��QdR駏ӛܣL��6/N�Z�/����U���:`,��'g���e.��(��Q���#�lb�1�M-v�c�q�J�B��Ν��L5�Eؙ��x��Al��ޔ��i	Á{
�t��濼���Li��xuhH�Kj�H���I�;�bwO$��< ���'�]u�+�a�T�t�/�L7_Uٓ=*NhY-��ЗB�>]�Gd��\ϐ֢s��sE��X^n-�	����㏀g���:���v!���T�Ւ��uͰIU �W��O�|}�F�*�Q���fѯ��3�ҥS��)!*&���q;�=p��#��fo��7��{�07�܋q?���#s�SW�kzЎ2��%1�,|������j*-pW<)�H���[��$ƽ�_��4l:7�4�0��T�Ǫ�c�~�S�Be��`.7���ً���v4�/Ž��ۇ-.��Z��6��wҟk��K40<�.�֨�r1��q��#��Ա����w.�Θ��|�c���o��9(�,����r�x��V��ib���Ǯ�w���ޚ���x� 9{Do$u�.0>eD��ώ�?�W�x\�Wq���]��&����(�2F��.%�Dq-�&�a�cۭhy3� �T�dG �1	���+�5b����5Ӱ򛱆��%�Wԓr�D�gE$��G����}�5��oDr��=%d}�dO|��qj��*'����J҆��x����eKk�����/ٟ�L�(h^�/�X������=�[p�I��#�Y�5��$5vNp_����Z{���r.�`h��-�KX�Q��U5�n	���4p�0Һ����}kt��;*�]����|��pPٜpޱ�����K���+�N�g!0۩D#��c�����@��~6W��B?�/��v{�&򝧕>�^�7��r_x0T�p�)�,��[�J�<%�ZK3vb�]6���v���{���M���ѡ�\{ w<�NJ���N.�o�i,~юE�j�$�CW�Z�����;,�8�7������oU���MK�w�䵿�3�*[ѱ�:;=֡W�`�%����.�+r=��t1�(�L:��Q8���Y&�X��$�d�2�-�}9z�JAv�7�t�ջ&�Z�-���Z��X�*]��#;#��ɽ�>�B��;�L�[Ġx4[I	ä��� W�v�@t�����g�k���e.h�p�g��i�+��(��cw8����/J!�Z 0P�ao�P@2���W��fD<��D��Ot�%��_i�Ka���E�L���=��F����>L������>�ɍM����l�z��*�m���I�P�>����k��h��9�����#��v��}ъ0#x%�'���?F�m�<�Tm�qFB�UՀ��e�iMzb-��VʇK6,�"�g���A"�%<�h�p���g1uޫ��NP�I7�F�u�7ӶEu��i��ә�^S��)���=���ۜ��G"�f[ؙ�i�Bu�h�f� ���^���t�"o�x9����:E�ٝ��6u�*�r�%��0���2d�ya�$!���v	�������N�jc,������O�Tœ�o���D����q� t7͑˭l�-�d7��PN=g�Wq�'w1�+���Sb�
�qu����sU�y%c�z<U��?m���������ͳ2T����7s��.�DP�
�+^�#@��Aȋ{g�J�`�]��l>4�[����W�����1jA�"~{ʰ/���g�m��� H&^��㱘jt���#؊��2�b��.+(�c�2`m��^��0�cv�^W��d0���?�%��ua�o����nO����+�Y �Щ��eg�\=�W�b�f���Ǘ�,�����ML_r�s��LL�^|�h�^T�u���nW�2'p���Ns���5��������Ԗ�p��H`.�g�s�I�oϥD�O��Ý.��'D#��m��_��`�ޟ�S���?Z���C���*����_����u�=`��g8��?��D��E8m)K �|/,v)�'��Ё%��qqɯzN��I/��;i9�K$�Y�����=̼����Z��+�(F�ݿ��5U
��I�㎧)K�y���HD��HůRy�4�k����N�-�c�\l��Q;ڣX�8����^���t/+/%�O/�ؗ�i_���-k��M*�<�柛w��V��:*J����6n��& �7l��Q%f�$<:v�l$�����/Z�^D���j}87;=)˭��[�4��(��tF��'��Pא�Rr�/�r���=d���n��4:��Ӌ�(�;��zAؼ
O�Y�0r@�o*84#�:oG��3~]�+���v?#%w��P��˶����mhz.S�0�D��=����:�^V��������%�Cw	����fI�=<�<�V^�qh�Pƍ�/�o��g�����T�+���nN�4���o1��l����zÝBw��΄% P:RԾ�Ƞ�"�u��UB�]>�[Wq�k���|���X�P,�����>��7��g~V���ggF��5AbcD@@%{��A�6"���OZ�e��m�܈���y�}�ռB'�������ʖvyR�y��	��t�'ˏ��7��lɖ����Ĺ�#�Tω�<2g^-���>䩞�۝b;�/�&���j���� n9:z��>�}Ab�\�o�"�):d]X������۲z�0*<&���mSIΚ����̄�iZ.�f$~�
��m&!M�>�xе0)�;�8��(t04Y���o|��w����7�c$17G�4��Wo��Ϡ�V_�O�r��I��&L�&����+�;:5@����-�����v���<����Y �\Ս酜fo����<j��Q�g<���a �3�v���l��M�l�@p��>��g�����u�ߙ��.�`��c_��X��	vGWu�*NYE(�5g�X5���!�����g%~qz1I���t~Q�}X2�gmmý���"��^Ai�v�(i�'������o+�$�d��"�+�O]�кu����ڱ������M��}���1�肥�0:�0U��w�����&��u���� �b/�&�H��5DxX+/g(��:ty�f�e��Is���e������������ZVNj�]�mn�lq�a�K�I�{�P�`�yO;^�4{�-,���6z�B�!��c7R��!�6%+U�����O�p�I?í����7�/�Mf0/%���):�@��	4Q�����F`��6q�-�ml?)��c� �Q���A���p�g6��$���
]��}�n��)�<N �^xzG�h�i�k<���9Z���g�;�9?�;��y(�>���5�C�����Z\|2g	I��Px�n^m�c��:O� �j}1�s�F'���cp��h� yؿ��S����;s����qI� x�R�0%��EԐ3��(�@�[�4�+��:Q�N@�{��6g�:��iQ֯RpVF�`Ʋ�l�����_��f�Rv��`���a,�2�0�JmU����9K�4w��B�W��5ϔ��=$��p�BLb���E�VBo�#���/m��.<Nѳ?��.~5��9=k���g�~��֌�Ӽ�I��a۽E/$"�l�W�h#����z�j|e"��m<�'���E;4��e�7#��|Ņ6l���+4�BuD�8Þ�+ę�"�gz�H�❆q�j:t���
x�S[ܕ�U;X�X.��V�WU�,d�:���E�a���	)�����)e���T(�a&>F�1!�y�R�PB���)�|N�s�h7Ȍ�s����D���<������QxK~�7.xV������H��[b�ou�����4q���>=�a��F��Uȵ�T�N��,��p8�b���ex�A��)�i��mQ�FG�M�'.��LaOJ�<�ļͪkb=W9zX���H���� �����-��ǳZ�����2Y:��d�bOդ���3�Fc������E�����D���W0�L�Xg(^s��7d,#�t	3*�/�K����ሺҧI���~����=$�Uy�n�K@x��0� Xb�j�z�>�G�-Gu��M�C�����fnc��y���L-Q��!����!�����u�"�I�׏/@��muk{B�[i�t �9.ӓ "���8ݨ���B���DbAoY��Y�;r��k繣�d-�+�X;I͈@��CA��=�O���C���.2<e�T)bJB�(,��i�Wĺ�/��k�0J�)��"^ >��|�-��S8��M5���Kk\v��1���_>�!|��^mBE�I|�ṞM�7s���Ck������EwK�џ�0g:X��^:�+�Q�2-�K������Jsv���|wFR�Q?-�ԷRN�5/��	R�ʰ|�
G���濰n?�1���������m
F�ɇX���$z@Y=r��Α�i���M�W�)�si��K�\���+?����+C(�0kΒ��v�Y��Y����S�����r�V{�b]t�����A�YQgE��3ot
Z=n��8S�$�����Ay���<h'��χ:�IE�lx`-���|�X��p��!f��������G���m�h��(����9���`��$�]"�������j3F��6;�����_j����Ӯ����'�/���('�68=�G`=�N��b�e/ t|r��|0�C{q�J������(e��N�]fg�+�����b@R�40!��N���<�l0$2�A��������tB�8�i�NR��U"z�'5K�kj�kX{톳�EP��;��J��!���~� pp������2�Kx�;ͧH	_���u9�T��TZ�.�3�g��AM����yӠ��(fȪ�����(�:���0n���n�q��_��yU�a'��{��:��@t"9�ǅ�����w} ��׹+������x�$��}��`�����;&�	8�gZ-h96_���j�eD ���F�E���6Xo;�7N^��&��57~:]7"ەF��3����� Sm�t��[�(|�=On]?�.�|Ԡd?�H׾��G��)�#�4}Qgr��&�Q�e�<UQ�?�RZ2��_����n
'F�\R+�����R����0�����Nvx�\k����h�0^L��,�(�.Dls��bV�E] -�ʧś�#܉Y�FFD�4�٠�W!et�6�v?�e\Sї՝>~x�)vJ/�Vi���Y_�8�xz&�G�N&�>�ٯ��l5W�>�����Ғ�9K6�����_�l8���U���u�y->{�v��P�x�+�:W<١�&� He����pU��̟x�"������G����n�>&�P0&��n렫����2�hp�/���}��y�k��T�>����;Z0o��l[��݇��(kq{]i���h�"}t�~����gA��Yn1�<��6�Z�EVPlV�ĥxNRZ8U�����C�z=`+����}���#���d?N���>h�@旟_k�k*����kV���G�;J
L�����ԩT�\��z���'l`��i<hzs������2�ݬ�Y`b�e�[=�C.'��^D��_-��6���u����f+~1X}Z�fl��y_=�z�%M�$�D�U(�I�L�p����J������=��j� Pm��;�	�s����g�_��l���e�%��c%\C�4�d�Y�I�}F���\��/��<+kI�[�������觓�����Ɏ������~v��$N0<�o��1&��i���������������#�DT��w��7E��z�˧����[ݕ8k����3��#�P�ˆ!I���=�+Qu�-��+�K l��j��D�7���Z�R�Q�W����v�TZe�|��"�͌��ۥ�/��j �Z�(��v�݅5�W�6�p��Rbh&A�U��_u�[L�-�d˾a��c�m��Y�9�p�
�'�����H���HO3�*Dq:�n#�@hq6��g��v-�s ����qW�'FN.,�C�d�R��Ϳ����&���L0��'Qa�����������my�prQ���T�[���~3v�!��2i�0lA�����M��h�5�
Y/�H<�M�i��>��d������K�P{6�c��h�4l�a��� ��,�����&#�0;�d/-���oLn���� �T.�
��)�e[?y�X��p7���+I�k��ZMt-�cʡ� [��c��1�	gR��Ϫ�a��rMP���Qi��?1��	�w��*ðׯz�'�f��[����,j�JI�LIl;�z߇t��-� aUx��ԍU��>���&" ��� ����Z`���,����vՇ��%Q����T 񖎏�'�-b.*<,UE��
�\�D�&�.�D�ِ[�����hdy%bF�"����~7  u��)/�����]'�K��><�)T�(2֤ge�c������F,��hښ?�u�p�|������%^E[I��#���;u;�ӑ'��~�F��޳�����dw�20�����:��Ԯ@[���oa�9W� g����g`K�_NߑT������u����R�B��
c���m��B����6n���m���*�Ϳ�bNۿ�At�!�R8�^:��lvO%�����}�,,�\�J�$>�[mu�KڛR�Khk�,���3�ծ���)�D������U�>��ȉ�/�̞=:�q#����&���`Τ�bq|Y�=̪�5�Y�9��E��ń�����r8C%Um���+c�bq�  X�G=��.��o�.����)�b���} W�h�0��l�\�Z�u��e��*�=d,ea���N{��g�7!e!���_	O���¶}�9���{�z�\��(���@����eE��_r'g8�R�2��	aO��l1OXP�ҕ�"J��Q� �R���e���X���Axh�^ÿҠ�Z*=�Y0�b8�w[@xI!�^B�+f��F�ui����(%/��k�PK[GF�_�8>�����K�	;g����l��;�+�pw-t@��5c�-v`r�)�V�ڽ��޹��Lr�X4U �oB�fY��3DJ��pH.�[ɬ!�r3'��u��=!��,���L��z��R	����`^�,�{8����#�W5���g{�����{3a���Y��Ĉw����w��F��F9�#��>��q�5DX�?:�R2̚���#�^��8�Ͷ73����A����l�M�]sq�� .�=��'6�_�1���82��P6�Y�I�t��L��.��fڕ�q��{+̩y�z�1�HH��s�q0���+&~V�'�w��ï�k�����33���@6��%��ul��
��r���=�h�� �!�Y�a;�Q�O�,��˰d�� �i�o.oLx��J�l8�2�*�g�L;%�~ì}�	\��u�OL�+#�1�������tħ�z	_ȥOY�ʀ�*�$�� ^�F�^���Hە�w$/�?��C�m���yМ5�PPQQъd:�Hg��A��W2��g��[�BX��.�7M�u��G�r��a�-K��6ԥ=�k�)�� �*�*vtIG�2b_��v����8�V�wZ�i��@��JWUc�;K͝^���ez#���m=�2�K�Ql}~%bOU7�!�8w�2c��+��Cz#��ۙD��2;�.^���3��N 4��4DC&�3���\��|��4'�8l&<$�>f,Eш�Q��'k@�Æ/r]��B�Q8�̧A����v�-��^��H6��X�!��RUt�5���0]%/b���)�KU#�ȧ�91ur���P��~m�P5���@a;KS�`�Ta��edo8��)m�
1� ^鳚7���f#|;������:��'Q���<c.�p��ɦ��O�5/h^��u���qP%�i�0�<%��R�T�<&+����eH1�J�߃�����̝��䇪\��z�~�
�S�e��@W\�wYRƨ�����39�7�	,PG���09���7R,�0��?>g�������j��qŊA��O�������zf��ay��Ō4��JlI)ϭ�H_���)	�11�s s ^T幹��p�2Bu���
K�@�XT�w%�?����r��u+ L�m�����]��C�W�MX���*��c7���NJk��@E�뉯(�]82D�1���c[���]��̃\�=����U����k���z�ׯ	^7r,����PԴI4;M�xvƁ,�~�ՙ|�_eF��N�w[;f��¯<>{����(^�_�+K�����\��L:�g�m�P�v�0c+����4d�,7�����Oosx�>;��M����39��|��:W<����U=/~���N�!���C�觤�$DQՐ��Y�w�C�І`;H���� �a.[�n�P��!	��	�!��b�X����NN��F�57�����N������YZ�"_��k���M�64�㭊�t��fE�s�- S��� ���H��a/�]����H\/���7�8�)
��c�f̺�pK�d����b�U�+�@�ALJ���=����Ioq�聛L�PҶ�$��%iUFQQ�>�T���X�#ϟ!�{>��	l++GQ����q
 �,�%����I��3���ͿO���I���q ���
9�S��*��&�Q��y�ÔLN=-r[��'���� ��pj0����mw�R�9���'���ڭ�VQOH�'g�`T|�*ӿBA�Б���� �?ː�:�;VI��A��s`��[;|J��<�Q3ʒ�ޛ�>����@�X!��r4jy!��!W�(��v���a9tݳ�E��;�]����8)��l8c�1I��<@�*�*�I5�c�F����y+w�~�R,�qK�(0ߴP�	����/���a�91Ǵ�:�GF���QsOA���&,5Nx��BD/	��X+�- 8n�[�Z����1��t�'�Ff�R�4��,D��j��7��K=�&��wxB�W�8�n�������C�K�V���\�}�Ȣ�Q'`f��縠�
B,+7<x���I:
:;���O�G��:�y#��p.+�t���ʥ�~P�Cާ�,.�K���W�7w��c� �8����S"ɩ9�Yx�]Ȥg?���Od�8��^�a�������*<p�W�>v��)4����m������0/JK
���,��z6��ύ���?1��2j�A�FG��҆M#u!cg�M,�
;�㷼�T�bw(�UZ�٦�nT%u_Z��v(��ܞca�dρ�?�Է�LW�g��6��&eN���<LG�5�eM	����7�(#sRR�*)*�y�&K��jH�Ff�%h���m�6X�s�6��fSJ��^��e/�Z��Ր���^����aj��[Юe�*+ϝ�[B+3}��,<��WwB��6Ub�_�2�O<IOcAPz��P]�Z�<'�0����j��LU�]��a%ۺ��gQ]���E�2S��v�	3��RC̸�_�(!Ɗ�z����b�o/3��D1�2��d�3�_s���"u8�f��;s�Q��7�bPw��i^�nR`�{��ﷳ|����/
z`��~���l���S�êV�;y�j��#�=g{��AwV�l�+~"�̈́S9�����|��&�L-�Xz���8��A���p.�y���0!��f m�W9F�R�LB���nH\�f~{
$��ma&������WB�g�k	(Z*U��	���|����1�j��]UyS��*�i��B6Y΍C���Ծ��x��h�S�z ���̵�#ۨn�J$�|�MA�� ��gu�Az��Z,l%�
�X�E��)}�)�k�W��ĝ���ލO��	e��p�U��c�'j4b��8��c1�uϾI�Z<��f��Y�C����4����]n��(_E����x5t�ʿ8�o�U�#Z�TX>�{�x&!�Ľ��c�?K�*P8%��ʋNV�$�BIڰ���?��lb�=���>f��!Դ�u1Rr�#������OjU��(�y�y`�ݡM��<{.�*��? �� �3q(�ϩ�ؔ�N̽�4���&x�O)�V����.��Wa7�h��S�R�+���
 �
�.�R=L��;ޅ�Px����_���p�=>��Uϵ^�Ck��"���|��Wx}y��R�s%��v�C�o��`C�yb��z�W�ae�wr��o�uܟ�۽EW�+{~�Qj_6�������<�0l���p%.U���[?��Br������q��¾d(�GWv3�����NA���n���s|T0d�˷�z��wc�ZC*%���(=�O�2sDy	��~�,1��O�X��xL-��j�*v	.�N��\R�#�^�VD/0g���S����i�f��|��8l�f+�D�����z���#�^:�$�O2�L���@�D����6��p>�X<�S���j����h"��be�@��@	�"�u�71��ka�ف���@('����WВ#�����PY������)p��(��M��N ��q�`����(t09j9�C�������2�	�
<mya��`�*暱'Gk�R��ڄ�4�T��V8[�����ӑ-־l�*q�{G
J ��QS�b�1@Z�R��@�ǫ�~⦉��A5,:Ց��]|9 ����Q�N���׫}���*x9�m�[����:`��33S��6�MS���ѐ�Z2n�gvc��-Nʝ����oK�D��J��u��&%���y��J���d�nd�^��x�=�ĥA@[ۋ�l�kPѴt�F���H�/����]݁�ɇNR��a΋�K����q*�|��՚��R�|���jP��2"����{J���Q�g����dr���q��-���C�s���:�)�z{@�( ��s�w
�4/{1�|��/�0R�:Y�nV�˵6�e�h�E���� ��C	�z3��K�ڵ�z9��f'��a(�t�����g���i�zh����s���/��~א�H������r��=��ZЍc�'qh�'���iUēK�ID���oM˼�]�A��1>��deȌ�����<ɏ%�L�Z
��0�0>���D�\%.���	��	dQ�>���I��zd�*ߋx��r �����#�`V��!���8x�@�q�f~��MU�-��Ϡ7΃"EV�+�Y|�o&N��l#�.��Q����89���OH�IJs)���$j�1̺b�
+�j�ډ�,{ ���������N����,�
��B"J�#���Lx����C�h
a�v"D��/E)�� �/�e�J�L��a�]�`.$�r.�$�3�{�v+�A�}Pp��۹-�t�w��МW9��0�x�/P��
��ɤ��5�2���'�i��F9O��N_4}�ē�A���;�Qu��HU*�Vc���c�Z�e;�8B%f�p�3��ՠ�zSF3��hpM�\�8qކ'��qg�S4o���t�/Q�P�Η$��ݳ����ϗRs��8B�$�|]���]q���K�_A�'��\�O�%#�J�GW;6�DB�w֜n��	���<�kG�X�K)��补7��C����Wh]�d��7N	��y9�b�#U���>�k�U�n�ãj<����	�Mj�eD>:B����FY��g����>�<�#\����DY��lь(WY,�S"�ojL\�$��@�>�㔯���l|Bvv[D�@|vT�_��G�.8DQ�5nZ3WQ�߳wg�遚Li�1 ���~ЖX=�&��Y��hw���rI���;*ȷ��.ᰱ��a��)>Y�|~R���Jv)�����t�Vad����\��.�������O��*g��}�Yf��>��D<T��,���iw��u�%��B�zD�nӅ�~�$���.��N|��(��'�Y���Y�X+ܮxbw
m-b�e]�kH����x����y$�&�E;6�:�6�;�M�����`�,����(�z�6֤c~^�G��l�N�dj�5��տNs�FiZJ��m>��6X��l�-�?�FR����f\����!@r��ܷ<b̬->��>�1O�$�����6�n�t�(�H~�2l�w�!h�r
Ά��
��$VZS�j���v���b�
:D>h��p�~L����P��s�.H���)��S&��:�`ɮ{
͋>��w� ~�Χ��kI�����~�?N]�1��������n^1�rmIē畡$��1?�b��5kA�b(�^!�[���oI����&�T��yN$�8��?o1vK=�xH�}2G���Lf�&Ć���M���ۗ��A�k���"�AI�����]���o�X��{}Ôp|X���(
�;�3�[�D�m�2�J {R^�9l���d5���=�VD�}���Ώ�`g��&*_M|�8E!ܲ�93����Fc���	�S�M���nGc��Hx9���4���T&��X������n��r]�ߒ(҈�;�ǟ��c7����#1)p��=��>�}��Cy���.G�ʰ��?[ّ.�?9�e�(?�Z0[�m���g�I��?�����Qe_�pbM�� 6\y�˃v�hD�-���+��(H������S���|�j��Y&�:����rv���;��{������&d�j��[��l&@$�(�*X���I�)'E@z�˚�������q��%��<�Y�,��"��ƻxc�p�cm�
ˉ�%vztD]Ŝm���b�v������;��]MB�E�� O$>r��`ː�;"�h��'�yH�nO��������y�ޫ�����i���b2��8�/�"��G��`c��������۵���k�q>HU��;�"D?3�@�-��*f,��ji$���a�����t�kH{U��F����=Drމ IQu��B��R���ZƢ�Թj�en��:�l�;��X,�eI�(k�i�e]�W`�&)�Ƴ�_$lfdE���&��Ѐ��\qj(��wV�5W�׎_�C8#;�Pa'x ��bi�=Δ\��Y>��֦8�.�[���yb̽xH��3��.rL��n����}<�t���'���C�&5.+�oAi�z�--�|^�Όx�Kۖb#����5�P �;^��N�?\��ީ,$I�Lg��k�O;�y�Ѻ�KLȷ%u׭�
�!\�y���s��M%dUا�cNDVR�8��n"����r3�WGý5�N���:�~~�N~�;�Pl8:�z���!�뷏�����W4Y���hK���� �C�X�pW�� �R���%d��y�|�E�&ў{����yFN}��0�j���CRG��zXOe����DR�����a�Q�vB����W��FX��ؚ����4��>�VIV?�1g�' kuȦ*�$�-��j���EIJ����P<�����'���@l�+蹙Gˀ����W:~Tς�z���.��/g�.�Z�'�u��5���Gj郻v*#*�0��D��I�~w��X�[0KOs��eK�E��Ϋg_����Āt=ے�p�ö��¶�]:9M��p�xߍ�%E� �����g[��A*�I��x{Ks�:�	BN���z���u_�;\��mި���u�pq���$"�hGU�{ʞ��6��h~�-�U69u��n��s�W:�|�>e����j�v�p�9���ջ�ae���>��+ē�Ѡ�/\�7�(�|�_9��#I��_�4�O�ê��異c�&Ȗ�I�m��~9�� ��a�j֕��->=	u�˕c\��S�^}�k�b��ʳ�9���'9�Ī�cۓ��kםq�d˨����.4��bV2m�<9T4It��	�'��L~���Ix��J���S@��]�����Ŏń�H�U>M�*���xz��{ȭ*�.��Yj2����C�g��`��0��(�͒٪k.�kO�yF����
ӱ�-ql
�Ķk �!�u�ѓ�'�9�����O�O9&��5�^�����l��՚4�%�E	3~�:����v��p�$U��?���z�:	{m�&��+�x����.��2"0��VN��H�q0c���K�?��d����\v�Yj���6's �-h�l~E�'����dI��AzU_ᦒ�x��Y����U�ȜpP<���K(�`Q�f &�b�O׊X����>dq[�}"n�x��Fe{tݗ+�4}����$m�
O��3z˿��X9���%�Q0 �|?}�c��[�D|��b��bձr_�>sYD�0�_����IQ dFei�R��$T˱;8؝�ֱ+�������i����)�|�*3mt�k¸����u��JA�51%�Zq_KR�C�Ħ/ʄ��Ap�Ǒb�����+k6X��q��%�S��?�se��c���*��i�ȓ1O�!����O���*SbX���W�^����b��dWnY4G��Ϫ�}��O��yD�m8���1���`jnu���ַ�_*G�=Pv���n�;W�9}��%e!�K/�s��iɂ�iv�G� ��ΐ�T��?$V�1�QɳNx̓�R���P�������β�P�}���RF2!��Y��袷
iGTu	��H���%ϕ4�}�e(p/��t(���,@Iֹ���#O�u��c�E	a!R�.��}-g����*䔰ջ����� �gSA ���kE.��GӴT�#L1�t�ﰟG5�Wv+_��]ܓ����q~�n@��,Ȅ��o�h�+?fI�9kJ�Nc����71�ĳZ�X_	��"�K� ��2_�%?r�8�qR�H0°{�����Ui�Ǟq�$�Mo�����y%,�tQ.��&�27KzI��`�i�M��H)�Y�gJpJѵ/�gŐ�����y��_[����,'	-�+�[/��a��%l3 ��<f�L��XuX����W�ۿ+�[>�_���J���::�cH+�����Nb�U�|���W�ǠQ``���b���Ą�������]�e.Ù��&��1�c9��!��?w�D����o��k�kܱ���ѹ�f�+�S�A���;>�����ǿ������l��6��a0i�f�t]�4F��ޑ�������~�#yK�%>Oft;��qBvUtf�C��Y��jmV�9�T�7h��0.�����>�H$�n��S�d0�&��h����*,x�g�.T���TD�O��[_�,��d\��p~�ػ؞11^$��z�X_�@������-��h�ƒ_�&��ת#�=G�ZKؿ;��N�dje:���X%��M2�YF ���||@�h��iWC+	�-$���;Q�0+�shR2�Ya�����1��T�>�B�i�Z�['�-Au�HUot�W[Ƌɵ����Ք ��;D�l��=PK��:&�����vM�s�&.D����MH!�+���6�&���)��ǈܿB�Ğ�D	���TBVb�6�Z�t�/,6Y�%7;��Q���<�Ę"����fU]�]��L��m31�P5a`W �c�Q<j53w���8Z,NV@ҪXj�g�|�l�]���_9�y������\zT��羣c��0̊N�f��=�\:�����&� \�~�{��U?K��`� �c�u�S�{�T���w���u�J�k���R�B�|Y��}.��j,�~������y0Q�&x*�Tnƨd$�cLC�Џ&fK�9��`����_���f�G~��!�S��0?+9����W��
,j���i�X�Ќ���\�Sڰ^<�.y�|��D(�l��`�^ޠ6FB�ɲ�WU�%��y�C��DU���z6ڿ�LHD�ݏz�#y�&}2���)��'J��w��L
���v�Ct<@�.���fI�g�'R�)�,��9���d���}=�R�P�li��і'�VW'R � ��=m[�n�SuU.�,|i�4B5�����POw�*���A�Xh=�@7zGJ%��g��X��;�c$���X�u��]�wac	�48k�uG?O�/]*��I��Ug�2}k��>��E���i������"�ܲ�K��"���`�z+۝㻌���{���&8_�����lͿ���^��>��+n���	2�Ku|�wQH�'ŵL�q?ۊ�s��W�d
�gĹá���9��zX8ݤL�&I���3��A[�E؃���M�| A�Z(���0���@�nO�n���|K���^8*G���5�1F��:}w!F�I�1'o����Ԝp��>ԇ
��"S4����mﯤS�������.w�gm�
	�����H��9l}��]co@v��d]~q@����Ӧ��PB�������ې]�<�8!�����ªMAj�ҁ���|u���@�5\�H7�m?�w]��ɰKRwo���"�5���!���B�8t�7����d�C*��1�]1�'ȟ2o��R��s6��գ��� a��7�3�O!�Q����յ�lVY�u�@>=���Sm0w���,iDGZ�uKF��S�alH�g�	�\�Y#��t)i##��װ|>tQ�%���.���*wƺ�vL$������S��S}��J��|O�l6�խ:R9������z&�:LA�d�o/���<�-U�K��f��3����c*u�PO1�� �zH�)��C�JP/�E��������n�Љ.2:�1(W*3D�=�Y/�LHצN�f\�nd��s���;8b@I�ڌx�AwM��fՀ|�1̃���v��+�B�)���Tn�5b�s�ɬH�0�BPuH�Z�.�����b��:w*��H8���ro��߄��L?�Ա��ԇ-N�΂vP'P��uo6=^��D�埼�sҏ8YEK��A����/�9%�X�9A\�����7�樂�W8bo���C�ֈ��gK:�&��g�"�xa>�v_~&;КS���,�m�
�&�LG��C.�r�E�;;�hI5���?O�Y��un��~l.�\�:���i�S˹A#�í�S�u�]�u��M9�w�~���zbdH�,?�O���?_1eT�S��Սztm�����P�S~����� I3����I�D����Uʶm�Qv����w���ι����k~j{��
m�A�r �˒]��k���?�&���f�x^Ai�n1��.�n�o�����K?���G�B��K!S��y|�m�YQN��0ZUv�R�+�2��A&=Ny��f��!���گW��P���Jqk�[�^}���a��z�����V9�P�[�w���$�{l:�ď*23��w��RL.�z�nh�ICbv%�|Q^zqOC�M��X
�H�;�U�n "+ �n�Y�v�m�΁Q�miO��(�K�	*�	�&����0u�ƙ��|`(���(xCW�� g\��"��Gb��;�]7��H������MF��)��-v�D�?�����ւ���Z��9�uJ�-!N��YP�� D�&��t�������X��ܰ�X+_��C<�pK{�&E
9`2<��9��T��ĚQ��-�����z���������5+ѫT�ۗ��k0���b�
��S�w0���ꏡ*�٠����?�Fm�V#%"gOt�d����PN4�v��?���n(nY�%�.kJ�Z��!��w��x��:����R�uƁ�����w(-�5�>�$��U|�����Ј���� }$��ށ�c|�o-6X�l�:l�?Y����v��^�z���as�L��Q�e�o ;�fZZ�O	�{�z"$�!\�!G��~@MgN�u�%�1gi@dU��!s룕?�ᷬY�Kv1��$�24��rժ��h��}Z�P��R)�G�S PH"��9uK8p�L��y�!k��i$�F�Yʄ0���q`�Q��b����U^��+`ƾ	��Y�͊T��&�ϕ�.W��F�(�oG
