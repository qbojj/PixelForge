��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��Ί/���\�:��j�gx]!�q�C�鞪�ưk��<�t��6���HV~��O_3�O4i `�����c�w^�@��5KB<6���a˒:80p�Q:<R�4���v�p���$�-�WQ[����@�(�����=0�e�4���w2��ǁ~c�f:+S�cqUK8�E�������*�3a-ٚ����ie�k��T��`��#�/k�z��A���2AF�0�����b_Sw��k�֍k��pO҉Q��5�3o��0�t�%��J*��g|bzwnP�c<����nK��E]�I��)BѣU7"���<"����"�_k��}���Tw$��l\��m[��ʿa���9R??q{���uR������G�E��o��?+�������E���DX�����EQ["���3>$��+�B�wO��GAճ���eV�m,u�]pd��͛вݢr>����mr��z���K^������M%*�l�(F���|��ƽ��͇e���E�^�;%:�{F-i�Q�wM�	-����J�=H��*:g&+~��n��#�k���lG���B� ��.s���2�jIϞ�DN>������l�ҁ��N��3��(��v�{��؇�aBl�6���N~i�λB=C/�e��*>�"�R��Ɍ�88P>NKߙ������nh�[������Q��+oQb�S�d���P4���$%�O�bN_E�<K��8���2p\�Q'/�N|���d��{l�Սu�ISG�%1W22��`�},;ߒ�z��t8C	و�H��%�����j��J����S�8������@)��U���Li��-%�K��;5��N�����%�a��))[X�uL.g���Q�Ħ�qN��K�k�!!�R}-��u��o����vQ�&�K��<G2��){/9F�O>j#�Aր�/j�O��qҩ@>?��]i�y�֒�9Ǵ���3�c����V�E�q'N���NU�ANN�f:�j�_c��TA%y�b�!�g�ܥ�TY��G������6�����4�D��T�h�?�X��#󭂴D����Ċ���I]`����sg��0qO^��g�V�������+�0��9$k��&9��9���a�ݾa�fMܮ��N;�������*
��6� 8�RTB�\�4ƻ
����f2���Hܳ΁�	�4��dP��feϯ�JZw��ʄ/Z�vRM�c����\��!Zh!i�40@�Ȅ�H��揄_55��D/)��@�Jc*E6Į�I�w^�#/ۮ��B���'�¹��D�P�����j5������t5���G0Kp�D��r�b�P3xkb�a�� /!�����<��N��Y!R7C,�������#��4g06��������s<z����H�bf���7�`���� z��kxb���]�pg�%�[M�tr�D�ў*�W��l!��܉jѧT�G�A�\:z��hw���ft�`,�[=�M�*-YO���σ_�$Z��a�!έv�VlIEj(�1~"b%q�;�=ص>��>b�W�RI�:�����
2�\����LY&Q��]�S㈡�ȀC���ɏ�v�_bE�v#���Oq���,�#�͟��誃�`"�08��K���JQ"ռ���}��O���8K���Ԫҕ
T�³���b1�z�av��֝2j��L�|��>�4�v�;���Fax�.�8�I=���@Z��5o�О�<A��H���3���s��
��%�8�0��"e�\&�u[����i�Tyu:��|�͎k���^���lg7��e���nZxk2�=��C���uĔ�!��M����3�O���)�`��x\E��_�%c��+�A_��� `��������Z�`�Prb�^��f�ۗ�g�hQ��G�Uŏ��wӝ�mGU~2��/!�q9=�X��w��D���T�	������XD�b�j�ɥG�zL�'�}v\H��&�8�{Ӯ��*����/�n6Hr��Vl���n�L�w���u����"�%�C�=� JF*�XJ	L
����UQ���+�56�hL��ݚ[<�ɗQ�q�cJ����R+�Zj�i�B,�Zb��wx������WR�=S��Y�x>���+ޞ>C
�R�����^]84�Rv�QcLM����ffF]��L	gs�K<�h?��/�"�1�`�H�׏�U�� X	�!P�<|�u���u�H�:�P)��>ڒpnh�;�,J.ۡ%sEJ���[��)�a�P|��tX-��_N�V�
:T�˛���1.f��Ĵ̶o�m��$���O�-{M�\�J�.��xm*.:P�� vj�4!��P��.��[LT;����e��.څwjt? �����8��(q��GQ�뮼:�EŔ؂U����W���q�H��t
Mj&Ҝ�W�� �J�]?�D�Ғ�v�)|D�\����!Sm�$b�_ֳ�% (T�t������)K	�	���7����gK�Z���2do]y3�{=q���=HOU"���������MTb�qN�l����:����%���P��p�����]����gݮ)a����%��d��"x�T+�&*UD��Hݞ�#����"��~��,�*���u�C�z�@]K}���mdr^����?-MJ�W"�gx�[w�k {��$�p7��J̔h��0����ăD�t�<�>b'�:��o�,vF��埿���	ך��MF�򽎷�E��Ӵ�(}��$'���Go���+�����W���(��i9�⃤�mϽWJ�A�N�n��^|���c��!����7d��� �����);�y�>pLm�� �0N4�����"�"է	�F���V�����(ᴙ�;�bYaw �$ D�BN�o�3��IG�N�ٟ�%F��T�X�g0:0���k�D��[0���
1
�峫���%��/�t����I�ܹ�q���U��P�?�Ml�D�J�.IK�;6,4�9�k�B{����+~gc��g��C��x+�(�,��v�c@$����X��E��b퇦�QwPg)���3_�\�1%�����1Y�I�K�}��Cc�`L8Z-
��#\۪�`���Xe��~g4~Q����~w"~�;0M�X�H4���՚I�t���ǹ+k��w��(3ّ<���L75�����S�L��;�;�h�3E@�Pqm�$T�����-�.*e�<��z8�sU� g�@���	h�$׮+K�Ֆ���� �j��\ވ[S4���tǚR�o��(��m.cF��l��؈zW��+�D�#3��g5ɣ��6�G��4�����dW�,� ��YA��-Л���ؘ��r�kW%�H1�7U{��fݐe�:�&�Yv���w_����vѲL��:B��)��(I�;/*SH:��
�0[�|����$����u��l
R� ۉ��Y_��8|zY�1㷖{Ɵ���Q��IH�T�8�����C#X+�kK���3�/�����Q�=� �KQb*�s�<P�]�,�t����DQ'�dr�;a��t_�x�T��x�[�/E�`_��u�8��B�:��S#K�O���W�U�W�J��GЍ j�5ۼ���R)�D�)5lo�/ڷs��k�+�@\]\|�xc�+�`@ap�|hpM��P�2]��!��!k�߶�B�A�@�9;��6'��Q��a�0��'���d�`�@���E�;?Ғ�j��%�.���D��x`S���}��]���3��
���_�S���R��}!�h���Cƾ��V\~�ǒs���P���%i|�]cs���4���ؾcK1�
^�!����z�ɲ��\��Y�ȟ�U]2rK�F}���Ց�w��8
�NG��� ��+>/f�,�I��\�1j�l�i"L���]�$�I�+2�]b�ԛ��>�n�~-���@��?���6�	*	��U�yA��6O���KN���������|j�D�/�.��G�R�O2�Of�������D��1>�Z=�߬c�3�r���hi-a7�8֏2�Fx�ŝ�V"�]���S��P���Z�ij�6�v]�������j���8_H��ޫ�$����w�bQ`��2[��Z|����Zz/-�@&`!���-s�&yr�$���18m:�q��A�U��?���Dq���\Ox�4Um�\2��HM����ii*p��ɳ+R�7�[�\.J8v��5�6�x�9��Ď��ȱ�";ՇYf��sʈ�1eN�A9mҴ��c�'/��fа�VC���ہR��%Hq����eh��;g-��� q�Z����D[��ǫo@�k�J~��'.�	?&��c ������(-��(���O�Y�7��[w 4�r�|ԧ�7	��|r�1��>��4؜�
C�#�i:�6���%7��ٔ7h#3�=pԨJXGF6����н��+w����h��0j^V1N��/���=��Z�R1��������r}�C\�_��$sZ�C�y�#=�Dg�6��V0�y�5�R��^��1��A8��9�؋*�W��
�M�Ε8���}F��G{	䦙�W�o ƕ9�8�a�M���8?��������g����SF��y($2]���yڵ,"�$�Nfa*�'�Z{9��(���R!�0X�[
� p0��;4m�'��6���eO=B���嘨��`xc�����x�?B�7���ԙ�	��5W3-z��<7{����W�=���޹�U3��:�ޤVX�� ��7fz�~��<�I�����]$gL"�;Q*�޿ه��>=�t�K��8I���^S��l�߅}��{����꺱$
Crd�����pu��@2Wbp��/Bޕ�Fv#��o#��e�%�@5���@j�����J�.���V>�L��K'Na��a݁�C�"�qֻt�7��S>�S˝>B0U�lA��l�q[zA��]ܭ'�5��0��xO��3x2��Ҵ�/q tZ(��X�Dn���T�\&�Cq���'̗�׏5s��e���c!ΜQ�EX���m^�MM� ���m[/�QA90,Ț�1�G�$cќ(�*�&3�@O9Pk�;�Q�F�ɨ��i�y}d"�t0������?o�+a��X�;3(����Ќ�A�ф�	�E1"��v	�Z&�ӰT�>����%L��zu��?*!�Ԍ��N%�Qq؛��E�=�&
�<4.����f�ͪI��[�'�G��_Ip�5�B�n�>�	�=<�8�CUEk�i�2{܍�v�t]��_>�x_w�C�ϙ�D�G��(@�?Rx���N��K����.Qi�a�Y\��,��M�Qi��rG&���� �~��l�f�
�p}	}z�zAOA�a��#�*���,-���8���C����؈+�d������r�� ��`��K2�i��,�2
C�~s+�9As}����z�)H�t����.��,�f�j��^9���QW[>��1�4\�t�|�P��׫Q�B�"h� ��R��p�ԱJ�>R�����ɟ�>�����/扌.���x��O�b���,�hn��C{k�%ӆ�E�)CQm8�C��ivw�tf=D��fmJ�{��:�̣�c���=���e��ǸV�71���%&�4�6�;� e$��$�}�d��"|�_����G�M�Npvr����wX���ϛu�b��i�o�6VB��f>���_E3I�#vf��1`�Ȗ){ړ��Zn�nOv��s��]�f**�����j\��۽j�,�o$�(S��ҠV�&�ܪ@�
���bAy(�n�3}��C�m��F+��.�� �QE
��#�[��2�f�)͍<�vdS��tx����l���ҩ����/���c���E�
J��S��xۭ@��.M���|�h����f֣�	l��m��Dr�`�t+D.��x&���y��ː:�e��61�"J�Is&����k�T��\"8b�̬��5�g:�����PJ	υ�,�2��Ϸ��f������|���5i�lF�ͧ���t�Tk��xؘGd��0E��m*��=,%�W{Xk�z�#�� ���#M�X�xp�m�`�^�J�}�/�הX(���8]�~�X�g/�0�{8�����Wm�^�~����z�?[R�;q��CY�	�9�꿳�"���(8?�'�������T�� R�k��T ع-sl�T7������~1E*�i������w����ҿ�O���J�/�qkB<t'�m�e��ɻ���RRD͝tEw�R1���)ԹA�0�G;�����qS���Z�I�l�!����G��p��˨А	S\	��ZhC�k,f�$��,����N�V����H߁c�f] �vQ-����6\ǝ��S�F_��!�m�A&y�0U\�,�ƞ�pH�Wx���B쵗F�Li�� �(���[�U����196�ʹ���>��We$T�j��jm;��؂&�z4!�W�ϸ|@��<�"f<_��755�n��Ǿ�Y��H�vj�<���X�I��|�3t����x��c�Q��!Z�~�2�P �S�	c4�ʫ�[�E�q�_N�s����@ݼ�~����^h`%����,C[XL0�R��kܠe�	�i�Sc�{[H��UQ�-|�)n2�L��Q��M}?����F�AG�c+i��'$��h�}+�h���؄Ͷ�-�ނ���}�c����
N傋ǈ��-j�e,s����.]m��M��'�� �IZ:#�Å�i8<3Eq}Mf푾x�ڇ��P��/�=���H�\p���.zT�G:nު� �`K� H9�Q1��J��x�Ƒ���Ϙ'4�e�:��-���+�Wh���֐o�0�n�M�9b#3��1�l{"�
$���;�
�e�y��!�v6�8uO���rM�����ѿ~�l��Cﹶ�>P_��kWy4mNҝ%���#������P)��b�X����23�uH�8'1(B�]&�6���5��俌����*�^����^����	<o�/�.#�MMz"<=��W�����z
�c�:K�H�	��֬)�lp�V�|�0#� ��T��No��>[�X�`;�C���Df�;��:� �8�N&#g��s1|��y��9�nU?[)�\��ބf*.����\au�R�$���ܺ�~� �$뫽'; i5�o���G����O:7ƫ�(�X,kK�X����T�f���R�(��)'��m�M�&�U�?GkO�e�IMA	�yƶ��y~��7���]6wz����8���M^|�i���A� �C�M���b��{`�-����4��8l�������3F�PH�v��A��W�թ��ˀ�4���ͣg =��l�\e��O�>Z�?�2֧iF����B��q~�L���,.⳴���ļ�<���ɐŧ�R����M'A�[��̷��[���*.5�X�etr����R�&�HZ����#'��݌�l�@�pi�q����{5�F���_��	�{�ܤ�x|ld<Ą��)��b��c�~��9�Ƀ#��t����bT��G˅��@��i<�ș�/s�o`p�= ��Le�v�,(��g� 0����[���/R�ܟ(Ǘ��=Z��cmS(��H�i�9��m7U�����{)���̹��$��x��h��W���'�^z^Ej��	C����^m��5�#]=S:<M^OF��ғ�w�Wm��nBG�є��^ʢ�e1�w�*����.�N�;{����0mX�)�qFS��Oy9Zõ���g��&�7�8�%�Hx�>��*G|�k�r�2m�?��԰�Z6��sT�+(=�z�ǻY۴�si���{��C�+�C���,qOB�ʎ��t]��a�ܕ���4�{P}<�	eˎ��=q-��ݭlz�+5���Ӹ�h�W��h����5���9�@��jƺ�.�;��ǻ�\a�7wG�&r��"�c�#�Q��|w��m�B�V�-c���+l߽Fx*�� ���G��ʴm�]�ڪ}k«�E�-��]�-)XjF�����c�Ը�D	�:����D͘Ͽ��*��&��	u
~�́�V��!�!�L�k
�:8h c���|]�m1� ǜ��'�w2��oQ6!���T`�����羁�"0��{^��EU�,�Q檒� h�,6}��V̺s�y%ϒv�>8k)l쇧�P`��M_r�)~�%Ŋ��;�p�_��\ڪE���؀��2I�p�Tn�PU=�H<g����;́!Y���'YC��g�	�{�k��܀�,�;F��l��v$���L�A|ߌ�S�!v�j��
,��~��U�"��BQ����'�VW��S�=�A_��v��~ Síb"�ړw��Ӊ�Z�0��mF�� :��DT�%�]�ˑ˟��n� ��#\#�v����no��Ւ<ƨ���υʁM���߂��j��oo�}���mI�.��"Vpd�|�ˬ%����
q���ǏH�tC��+���E�~��E��_�s� Ag�#��䵡��&�1��s���꯾?��R�PFS|��Q��f-[�N�JD�x!j���h"���}�'�d�|4>���9OgΪ�IU-y;x�Y�K��р��)�2����0��_�"?$�/0��r�J�4J�9��lO�8N�� ��^\1kjo�-%�<�2[��HsjN�$ ��c8����P28�?�
6�z�Q�������Xd�)D��h�%)�8k�f�h�,�m��ÁV�lw���[Y�;��1ڟ��i�UZ�E=�/�<B�值=X)9�̔��lX
ɮ�w�kȚ�N�k�+դ8�ǜe]��U���x���˲���ċ*��(=q�2��>����KUjF��S�.s`�G�Y�@g!�X�YN&�[E��9|0�z��Hd���ȡ�D.�8G����h��I���ୠ�8͇��&K�Ϭ���]w��F��h�1�J(E�<��a��N�	��*�#��\�[3�x�t�&q?C�k�m۷4|3%�.���!�p�
T \Q���E����j����:��q��ۅ�t��S�n�� �!�L�_����m�=����z����+:4�W��í�v��4�7��X���)��ȝ�A"�f��81B�N͕��[(����g!f	y�����Ƣ�U�P�%z@{����&�Z�q?����q�jon�Y�d�8���i�~fcL�v������e6>u�D�A[��jM%��N�h�S������y���܎"����eBu�i�v�^��Քt7��_*�4�6TA/m_�L�XH2�����%f�a���t���]>2��'x���|���{7�Q0��\8Ȣ@���z]�Į�q?��Y$L|�]]~�3n73����鸺����8[͟�9!���U�<k�SzN���8E���9�N��Q`�i����;���&`��6F,��Fh��K� ؋���AV���ͯ�3y ���4���� ��p��SP/gyT���G��[@�y2z�!*Lq\�Z���eN�qr��Y<_YO�����+��Z�<y;��9#�w��wp" й}�vc9���b8����3���Aa3sC���o䜐�;R�u~���x�Kr�BU3����aM5�Ѯ�^��#�K�N�h5���w	B_�}�#a��0�d��!<9m�T90��MU�v8���9x�ؠ�qbM���"�4����y�������� +/�Bn�j�#~6W��`6`J01��с������=R�h�3k�q��y���;���Bʲ`�/����%Z�8(��|�@ �2����6�y5h�I�v�\t��EJfz�pj�a���c��:�@�L�M�-N���,�q�c5��������(n��o=[���٣'��cI��^b�Y[�`Րg�a����Tpͳ����]T�2��r;��5�����K=��6������Q�ث�F�t��+�oz�0�4�n����ds����QO�����w[�D��t��
�aC�L�R���N��G�p��=䍝��MȮ��{���{h҇������}�����T��1!�*��!5��~��^�]�j
mZ��P� �V;�v�R���OB���0�*�lb��A��Z/<������B�*�%MqL`�S�
��M�CS�21[�}o:��Y1��0���W�CS2{/���:����{Q$މ�G���?��l�*���UN�����J�*"=Ȱ$�e�!��L�{�z��mS��e��V|cJɌ�k���uK���̮�Ç���ȝ���b{@����,��>���y��>�Q��7�(�""�m=��Qd>�#����B_<����
��~<���spr�E���p��Rf��O���he��#��B.kÎd�D��]Lӟ�����zW�g��Q�[�pc��.�Nk�2I.sK��9�Nv���C�;� �'�Q�\��6'@�:#���j��U9�߁�\�$}����F�O8'�;1>�`�d����fA�%�fh�wd�Q�<�.�:Sȩ��
kg�@������*�9VV'�����G��@X�w0����K+�M$H��=���i}0�K���TXԷ�'Q����0�RehG#	�J:�~�]��*��l���o,�����*#��T�W�g�.=}$��HW���;�gyàD��t��.f��Aڍ�^�
Ŕ��>���6��\̣�ACB^c9b�keE ��]���N��iܤ���i�jqr��Pw O�8^��B��sH��Z�����P�ɥ�gN�6^��3B����9�j��s?l�4p��xf^�p tl����>����~���e8�8�([�0�"^q>	�p�����H���@������(?����쵦�T�+�P���)i2�n))Bx#1 ��|
�:�:����yO���r� Ё�:�� �cV��k���N�BD)i�Px�|"2�a�oe|�,	��c�q���%���zۃh��E��<,��C��G0�݄�L�?�+�1@-�{�Y��ʬ7<:U{'���M.7Ђ@N�_a�}v�@Af�nEˆ�Hk�ڗ�����ΎA�$;�Թ�]8F����3$�,�&�8�(Қ�2[█�۝0r\���]�N+nB��6��&�d�?<�o����@d"�	���ݣ8�r�f���#�����wV�R>��g����B�����_�ǦM`�3��ù�����$D�/����
}O�7"k*�Q�i��v���exx����C~�3�"�Z�j)~�Zh�#+�V���!nrxkѾoU����-MA�,��}
%�5���b����
'�+�[1���{��ȥ�~t5`d���/^�v�4WW���yHK��+�~X.X���	��WCA�������,=(83'��2�(���˽٥��rggVWz�(=�*0���.�����ǚC�[�b�zYF_5����%ä�����{��o����c`5/�lR�2����_����r.���F&���l�C^�B7b�Y� �@�#yu����a�n��n@�A&MUTgK�>���Q��������~L����2�����oz�(V��x
��n�Cm��7�_47$Q+�g�F�+��U���EH�hTG����y��TTT��J��,�Ƞd,� X�Vl��nQ��s�k�l�m~5Z����c�� ��3/!���	�\_n���`P8Ч�t�}W階j��S�5��\�#W:�F��p՘���������2�&�`�*_J2�3^��G���;]n�e5���s�X�T��F/�B_$����S�1Z�W(���6��0��2~�=�b{D�[�!���98yZM&0M���N��&��}��j��$G2KwT.��g���>�Wg_Z��$ �I��s�F8���yelɤF�c3����D8�ڴ!��VT��?�G1��!��^���.�u\'H兮P���I�.��D�V7�A�ܖk3і���`I)��)�(���ݘ�=�z�f��hUނG��Xh������;�0����6Y-DTT����'-'���m�@o;��q��[����5->�䠊9�YyxuH���e�$�����U�>���P�i����-|�� ��!����w�V�a���j
*4�h�4�P?a���"���G��Dp7�CO����ř7>D����x�1�3��\Ɔ���_� G�(��GD\5Hs �3�����M���=������0���O�~�G �1A?���NK��� 8(��0���,$Ы������P�_Wܾr�c��~��;��$�Ӯ���d�w�u�M&��m78�/��Y��7�m%D2Q��d� y����σ8���"B[�D*�G��ѹ�i@D#�`v:m�b>�,�p�8M�b��o��(T�ج.��c�Z�!��DK)�,]2�H�?ƾt�<�)�9�Y\hc�P_��Q��ay��7��B:Eڗ��̒8�Wh��\��j����&8s[�+��:�Sf�iE�2�۠
�Oޥ�$�Юb��H}������2�(B���>���hW.JO��B���2��@`J:�|ä�Q�>�ad�'��
z������Laiv|z����c ���#�����(<B:^hh	�1OV/���	�
�M�tD��{��$�q���x�C�����(�Um�~�9�#cٽK�*/e����� �$�{��[���k��p?�������GG�d8V_dY�$���F"����W���h廒�=������¸K2ޡ[��>MXʺĴ� ��*�q����M�(��M�O���Fmn 9�l]��^����U!c�,���@�Jҫ����s�W���N����VCr�0cޔ+kϠ�nQ���qI��|�H
�:�����d��ǵ٪z�GU�QqQNQl�W�g'�d��K�|�7�}���}؈�u���S�Bt�0��2pH}��Q2֨H�����(��=�0s��O�!}����1��]�s���[��Y.x�vVr�>�n�*=M@���lE,�SZ����E7`ĝ_2�*d�ݰ9R�إ�	����Š�9�{1��L穻G~N��o���h���p��P��]ڕA�AY��=�M\����A���W���ݯ��qH����8?]�gIHk�P�P<˩�OT�>��y�ÄLa��D�P�Z�8���'�?E�M���;,\�j�q��ї�}�1��G�/b�%�SW�̫B�M{�V[ɨ�P'�na�~�_��Ic~���Z��uN��#d��Y�
�f��mvPu� �:I�p������!!��~v܌7�EY\΋���.���I�d��^K%���a��-��Am!	,�&���N������w��U$��}�F_[�ߠ�:~`�|��V�Pax�-7��4e�vi�c����&��|]����z/��%��ʹ"ۼo�u�:0%�P�k�ȵ ��4|~�q�J/e^�fXUL�v\|ƉQ��z�7_�ȳOCgoR�X�?�y&v�U$�ݲ�:�$�#G>y=�K����ò�[��W�{ٕ������� ��\�VgB�D��0��H`a��u�z꯱���)2X�]
PK䙷��[�o�����'fխ�mo���� ��K�P�����K9su�ɔ`�'�� �m�+�LJ��Qh©m�\����|���Y���H�,8��^Z���ҳ�uv8�W'��A�2/��3����:�������Ғ�n���n(�k�m�s,[�<�B��s�2Y�2×��j^�c��}t:��-�(�n�Gh[�������2���g,��:E�sj壤n�x<�ƨ|�����ܕ1<�ʐH#Ū4f��i�P 7K���p�T�Y�5ܔ�h���K���a�!mx؟�Q�����x�=�v���-�\htF��I4�>�Ju�Q�_����/�S֛��Ȗ})s왷;N�ֽ((���@�4ԓ�c^�[�❍p�sJ����qB@�Ѭ����I����3������k�@�ӭ}��]*����L�4:�o�_�H�km���w�!wO��s0�@,���%��a����i���� 8�	�³��'��8��i
�����=ᗹ4�C]%���3QRt��y���.�-W�ɏ݆�{X+�?jTIq��Q6�b��'�Ey��.1BA���T	�.'�AŻ�|GF�PK�䭶����Iд|��^nȹ}�(,���h\�Q����ް}�?�i��1[��� �@�נ~���%?[Hʹ�2_:-����p�ئ��`Fn-4 ��|�hI��Ċ�n��z��(��ק���L�c#����OG��s�V�tϢ��=
x�!�����j�0vG��ZrճęS���>B��ɶ�S��v�Ba��0�Y�J�*k��������~�s��À�q�H�����~���㎴�P�`V�>�K�R=��D��W048 ���Dq���{�)�7/�CR�vFÿ@d�����x���	��k��:ye�|^����8�	@�������x�!��ۼ�%h�f})�꿙��f���
����܏�W�i�c�����RB��L�>F�H{���Q���;�I��e�|��i��ԝ�⃤n �	ڂ��TA*����֐7V��siB����q��AK�^����Xw�OVC�l��Ӓ���}�=Ċ�����
�"}�Lt�"�GSr/�����CsR�t7��h2)��-��w��7	VeV�`�a�Άh���n(]Ƣ�\܋�i1��%>�o�ցf�P�#��Q�w϶����-��+�~�7.���(0�\jp����o�1dW�!+w���?)Q�ݯR�����So���Q��n%��yAdJ	��[��P�$��Z2B����
�J�o?Y^�q�1�bW�m�*m��Xly�i��R�W:��AB��Y���.�������pM)���YM+15�!<a.��:��`M4����"�s�]){J��{�JV�t�x�;���ϊ?�<�>�-l��s��B����6t�{YҊ�n�5D%��Nfia�V	'K��u�Oe&(��1h<�;9�l}pr�G��@ �?�?Y�Y��GZ�J��H$���@�9	�7�$�����t�z����ƴ$�xtrvT���O��	Gd�?L�O��o��2�#��0w�@�����N��֐-�z���N�>�e�9�օ9M��#���������!������6�jmL(������׳�j��������@�X���][��`ǭ��EY�c�ܜ�Tzm;��f|��G-��ѕ44B5��fDSX&i�@?�r��A���Cd�t+#q<�G�U��F��h$ֆ��N}J�Ѵy�Ӓ�˒�_A�[�XZ߄�v���ɿ 5�39�`�Hp@-���܈"�Z�}�ƭ.��UL���
[W���l4X��7�<�����G� �˘1���s���]��'�j�Z#Y����:z�*<p��מ�by�#p
��[�� �rT��6��F��)�E6�e%a:4n41B��0��si�N�5�����e���Q��,�%M��&iT�p��H�%!	�9q{�V��߆l ��yy*��ӈ���N�D��f�؜�(�����������G��4x���s0ҝ�t}���"�&�,��v���3P���i���^+'hώYqʔZ+!H�/D����p��ղ���Y���v�BVG�a���^���=��H*ƫ;&	�zp�;�,#O6D���'J��uk�.�q�����}��.�c��l� yt��n�T
��%0�y�ȡ���ct����w[�8"U�I}YZB�e��f�Od����]�Bx���q��G�OV��s=)�� 	<���)q`�~M.���)�w_y%#69�R�[p�C���-P��W�~��_���s�M�M~/�MB]��{��H!������I�D.X�)���<�&�XZ��.��&X(��hlZ|���_4� VJ��_R��t���N�"�L�a�ժ�N`�
U`�U
�k"B>¿�'�ň=��B�^��
�{LA��~eK��u-����!~���D�0�z� {��C]{��G�%@;\�EM�#l�.�>NkQ?[
�~D�ZIH��T�շ��u-dy�o�1	-�КH�~ڜ��\$^�)�
�O�y*�����YO���H�Ð�waR��?C���c����9�&����}*���w�t��mM�/V�1PL�\7��� ��^e(��@�f�~��Q�g�&�&����{�P�xG[Y�3{7l׷����P؝��W��q?�6������s\{Tap��$�Z�9��lw��\�C���G��IM�$�ĥ�c�c�h��m�O�u7:󵨻p�xD ,����\b}�֧iZwyG��?2��Z@�J4t�F���&��w�ˑR�_���,Z	�K10e g���4,?�«����R~��D�u�ģ�jֳZ��ك� ����x~���f�&���Gc}�萡��_v,����#M@��#�!e+��]{mT:(k߰W5��Ò'�tٶ���cJ�>����Cַ�)b�$�����]�ӈ�7����(pM�5YhG���	�'R>�S�6bT )Fd���O���n��ŏ[r������Ol3�V�̭�Z��<,*���Al���@���5���!%���=�l �۶�pkS3�@��X����k#$�C|�#��B�p�T-g�uO�-����6�km��=��Ei��[k�Ya�8��1�c�⪩����d�^ؚ��X��լ k�h
��!8����M�O��|i�niɣ.<����;�*�m�F��
��/윉Z�E5I葥-��n��Q	��+vEl��;=c�I���01��,'f1�qv�T�08�{&�He������S��J�~����X�)�{��|1R��b"r������Ɍ'�,Ǹd���'���1�@��L�Ɍ�_q�_�<�ywm0�c�Ga��B%�dG��
AyQ5ф����Y��w�뿹`}���9��ӵF�r�(Lk�Ƽu`s�"y�7�Kd�H_aT�����ٳP�Rzl�i%��n����M���t@o�s�s�X�'r%�ZIC�QE�c�!��L^8sY�&!ņ+VDt�l�r ����%K�Qɽ�-)�^�w$M���N1E�Dp���8K�(��B� ��w�=(��֛;U�5X ���&����L�LlYf�.����_>z�	N���v��e9du}�.;�O;���h�%��7E*��]W[z8�W��/k��ð_Tq�-�y����շ�m!	W�2f?��}��{����p�*X+�CTU�}���8m���8�z��]�R�&��E�����
},Q� =�9	�Ǳ�{�"k^<Ħ�l<%-�۶&�d�Y;����_'f|}�LR��N��p-nԢ�kk����䰭�Ϳ(�.�WX��e��?��lhAY�~��e�Q�%�}1pE6Q�/�����A6%)D��/�3�n��U �8s�jZ/�Z�SĘ�̺��TK�~e�ՉA@5xygGp���;�Yi�ş�
޴tb�E�:�*⷗�0�s	[�4���Y�櫔�f����L�;����P�#�8�����4�9��j��g#��R�v���+��Ub,�I��FTڀ�uN�La.�45��s�G�n��O'+K~͐r
��r��3wB�B��O�E?l��fg��|e����ّ���	�$���	��yTXk6�L}�脵�T^>��um";J���6=n�"ƏeY�N�_�uƻ����BY,�7O�N7��<L86z�誼{���O�U�a��J����}Ïco�.���@�W�b�-�ZM58>%��j��s ��%$cۺ��Ln��t�l����ԡ��"sr%X����I��z�7�kz,{��=\���'����aOk,��ɒD����U���Z��*+����K�2�\6��C=��WV�r���`�NK��w7�93�����A)W��:���R�b���ȣ;
˞�j�S��wD@�儙���V��о�F"��(8փ�ee4����:�_��rhd�s/t��
�׶~y�kN�j�{��nVި&�T�w@��Lr꽻���7>�*j�X{=��X$_F6�����$hWA�(�n�jH'�3����Z2�Z�Ϻ.u-�����C����(��
%�_�^*h�roov������u�X�M���)Pw��Р�F�����T�1[L"���y�������ɥ���a@"�`60ƅήʯa �X�S�J<\����E�f�`'d��"�Oh�A5~I�X������~D0����b=���<˝̶o�XzC��"�C�"wV��Bb���c���jhǻYk�Gzl��b���6��:1�M�2�R������Hۥ��yln�����9�S�3�fܱ[�fD-D��5�
\��R�3�e��x��ԣ��鏫_�+b�f
��(q���w�!Iy�� �8WA�n�����WWm�g琜*��Bs����c�Id��/�q���^�Cΰ�}D�vu�Vdo�b��Q ����H����,8�g�y#�f���H�i7�P��6���R���Ǝ޻隢�	�|8`��}��0 P�kXu�&�b��������+0�S?�����_'QP%�]���7�
�����7D�&7[B�0xe��$CG	�2������%v��Z�ǵ�c�Ǆ 9�S�V��M��d��Lz�L�99���w����׮OQ��PS�iQ�.��`\��2�"��Bv���s�����V`f�Է6�����(ZOJ[��"�QKH�SP͏_�b"l�k��V=����&6�~(MN��\C�qx�����'�ˑY��ȼ���jdp�
����x�,�J�Ȩ�Ձ 6uo؀a���vc�A�` �a@&�rx@�Ԟ�����l�t�H4d��Jt��ys!�!F�����zD�]��\���d�%Y���@�p��e��f�9SVi_�wy�p]F������W��_j|Jр,�u�.!�)UVڭ��:ɞ��<�5���2�ⶾ ��S2�]��e[1<���#��3�8/n��V�q��˓!��iZ���I��#Y�I�S��s�I�9����޼���fl�W'B���F���e�RD[o�&`#�G��O9�h�i!zn]Z;[��(m������X��wU�O
*�kbf�{������拁^�����Ԫ]�P�~s����Un�-%'��n��}�~$�"�{ҹ~��(@&Q����"-2��̻Wa����E�ܶ:���)�<�a�-� �#�;Ia�Qw��:;X@�[It�m��P��q�_6���rglK!˱���Ƀ��ݛ�el�I���X�7'0.N0+�H	i�j�\��N��9�,$ڷkoT2|'�D9t�q�h �')�&�G�CCP��E��G���$�_J( ����YK��_��u�e5+�W��q(�V�,E���4rX�}|��di�	6*.�����
,��!��  �����2��w��z� TR�+�vT�J�WL�%�ٵ5�_�n� =��˘$lOȉ37����<�����ɍ#o�4w��Ls�|(@�I�{����|>�����Cԥ�4�XѦ�ŊNg��D;�c ����~ړ�M[9��(��!�%L��l:
�_�p0��w�v��5ui=��jޥr���D���$�-:�`e�1��d
���?ꯉ�a`	Fc�k�{E�2�(JKӴP�G�����2��h��殦"a�9;���	��޴���u��#��P�v�N��s\�6�E2�챩(�a��ϱ��eF ��"&?�������fF��RӅg?r5
��e�<���ʨ1ZBg�=N���z��v�Ǭ���Pݢ�>čԜ�)h�66gt���`p�JQ`0�7>
�5��=��9�o~3�~�T鹧��ٔk��53��%�m[º���nh�e17 5�"Qj�dOǂ�c�ɝ��r�_!���H����c��3��_�,0���$C{����޽�z[� ��#�^��m�&\�s���~�y�zb̽z��6��<xӒ�c��w�I!!�c�'�r� �'@���Rt����Ѫ��ek��Z��C�����^Eޭ��//���}�5��X�a�޸����'��*��h�\(VwB��������>�)������I���.��=��,��tݹN� �'&�t��:u�o��ڗPǉT0R0c�r�F7���u
{�7\��=�i���zS��M{#�|?^'^�u#�eo-�~:�0WIH�P?��Ÿ���jf��=_�6架�/������j���ʑ��z�O&�~�4��N��{�5B����B/���D9{%���@�$r��cK98��ɴe�h&n��T�:"`�Ѷںk@���'ǈ�00o
wVʢhxw�'�8#�W��� �G�A�O	�|
�r`�s�L|̪��������vp�������m�V;�[��r�*�!ڕ/�z���c
jD&t'��j��Uj��|�k|4|��^=O��n�����$�	��]%A�b)�*���.��U�ZL�����"������U��`>|:0\�u	��7��j�[�Io�=q�d����|i-���lil~�Fg��]��⊴)&��4K�H�������_7DSˤQ|�����b�!�/R�޸�x��o�jU�u���<PP�vI�j����
�~!4簂jx�A�J�-oG������Y�����K���ԎAL�ٲm������p�~����+E3��� ��!v����-ߩV-X�$�4�}SL4�Zu�}+��Ǫ8	�/S�b}.l��)��2�k�M\�K�$�����'�4u�� `ܬ�S}ti��s!��u"FMo�����2� [Ieu�y`�">e��c�/���<�U�hS��5��E}������f�->z��RāL
Q���TT9�O�4Ϊ9���[�c�i3҃�P+�҉2��.�+�)9[m����6W�!��:�o,)^�*NU�$���lL�>��Ƿ}4S�2���P93������HG�ÙZHq�1�W!����>��Gϲ���bb͔�4��`ᗦ�t6�iL��{}о�0er:*aخ�y�Z���x%���C-Fb۩�Ԧ�^av��>��i�jg�S}��
�CK'��i�&�Wm�¼P���[kJ'�bM�T�
+8��|�YOi�<i���ܬ�R	�0��E�1M���W-H/ۮ��6=%��+dM����U�~ �Y�C�na���R��I9�[�mY��R�)���?B��X�x�����u�@�D��ʭ+��p�솫jn�;��w�Ȣ�0�G㘍�C�3A��S���À҂�f[u�]���W� ^�	�=��)D����|t�4�D���� X'J��ADk}����!�n��(�(xɶ�7�p2nm�Q��#��=/�awXLj�/M ��̵���}��������GM܍���~^+k�$��#}h>�m�EBd�^J�z���Wfǵ�mX���l�����'EZ|��6��K�-��e;J����E�t�m>D�q]�����x����ԉmK*��`\�'�J�RՀ�f��܎��K��؉T��ٶ���A%36�r��lr��Х���������V�z`�j���z���4��-��k��l��Z���%�[���k]�mAw0�>
�3��|�*��R�w��IyPÚ3�K���:?�,E �w�\C��Wn2Bz�Z6����a�����8�k�S�#�#����V��tQEo��Ѧ�j��'����?s����i�4p�u0?���ؑ����
��p���g�@{�~�s�S�~�l�}����}����;|����ւF++_,�j1��2���P) �ǹ�h���g"�U;p��_#�!�	�����.V�D��y���rq�D���L�/Lm���#7y�1,�wW'���>�����0Y�Ϣ�oh^�}��	-�s7�Ʋ;�Ɓz�Q��uW�@M(�ac샔%E�bS�`�J䬮2s�	�YGA��� =MJ��{�v1�2A 5�dU�]��)�z��#z/lԅ�k[fnx��I^5��xi��{mΐ3彙�����Vd金�����: �hF�J0�{B	ᔗ�,lN
�=1|@�V-f�1*x�ȗ���Ùj�K���H��c�z*X��&#pS���4D�� ��ܝ�*8Osr�	�2����\�_V�r!�z�\t$�YZm8}�� ,��6 �Pp��"'T��z8W�Ҩ��W�'?�7��P��,�3�=[����t�y�ޖ>*�I��,cm���;�\�&�����}!�H��(��#��R�Ы��Xإ�\�̩��5�:[�V�ȐY�R������|���6	�?�p��4�����O�d�7�UvL2�$N|�Mr�]@+<Z��W� 2d&`���7*2��l*#�asZb�]�V+/q��-�� >QZ��|��v�4�=F��
����O�φ���R�r��p՜a���R:��7����;��F��;�9\��	�.7������
��;$��O�@3>���R�$��߁iL��]Y���"�*0��v�{�e��'O�D�����"�����Y�F��闳w &��T�ʊ��2�+BC��^����v��T&�P�����zE��B��:,@�&�n�_��AR�n���4�g��V�o�F���J�Md�1��'B�ٶ��^��Zឃ�����~{�Bw �1qdb���{��7��-g�P��	�o�\�q�o
߂,��Wj��#�B�(�i�:Lr�e_1�NֹmI	+�`�PL�r"��F�a�2���sLq�di��w��.3���G�#T�5d���_@or�o�4������V�a��.�d:���\b8��H�H�l�-���7$��v�Շ�v������]O#?(��*���48��.2uH��BG{$�(����L�P�5�Xp�b��'��n�������/�I)�j��~��*]u����oo� Zw�fc!R����<�nDu�|�\��@Ɔr`i�/��E�n�܊�l�����R4B�
�f2��۾�w��Jt�����LS�L������=#�އ$G&��-dBs#{���!���&��MUW]��[�T���4T~^$j|y�����%�Y�������̫��Y�͊��#r�b��|�&�(��t��10�9O�?^�S��})���4r�M�r���1��V�^�N���/LP$.��̾����Yv�2=�L%+��XR)�*g/T��7���0�h��I����a[���9�R�)�'UE(�5����
7��K�F:L,��WJhG �Ģ��� P��w7�AHq�2��A������(x���r^q�6��.晗L���m�hY8����ޗp�N� �~2q�&�_�u:G�/�z�Q��u�mo!N9���I�χ��`��c�n��]���Olr�a9%��0Z�J���j���~�{���%bUQ&{��` ѧd�t�ս�;U7��2��!)](��8i��Ԩ=N��#ݲa�m�4��I�{����}!j5�p�&���j���:>
�s��u��ht!��LԿ!�@��w��K� ��n��Ƒ��_�l�Aw��Q3��eȁ@�
f�{c��0��^�a`sb&;Y�^��a����t��Iϣ&�ɴ�b7#�`��� �8	�S��*�Α�b$����MX�ʅq���FF�R�C��곂	D�s��S?�j)�!��v�l?�d�_��̴�[�u��Ud��3�!����0H�&�ڂ��|u
��mT��'�6�5�̪�/�\'2��q@N�F8����r�p�����w�K�1�����ae!2L߉�����Ho�ɰ}�N��盩�@G�� �Gg�����]�@[��H�i"1��k١�*����{S����#�Jv����J�|��9EHz����9A�4_P'~�U�[D������QoI�r��9��_mA��tSa�n$��@s�]���āl�0F'ط�ױ���*L�x�����S6 ��3�_�j�t���fZm���Ͼ(���L�(|�K((�K1_�����a�L���3�Q�d���<FÕ{_�հAH�*��)L�Iu�ss|���0^筐#q�g |y%J��4���-���#ذ��3OX��v{%E)��m�EYG�8�e�S��=ĢW�A�IAR
w�%*����O�	�%�����S2wm�7���۷��$����%� �,���	�M459�[�Ŧ�֏��W2����Z���ùeOz.�C�j����>����YfZ;	�+���� *<��L�����.cf�������߸�d�G �Xs�!���.�!��b?�<:�Z9$x<�O��ê�U�V���0�r����qb�&-���O�����:�@�Ÿ�S�#s����>�-�.myc���l.������J�d�H�w|�úUG2��G�k=m�I;)w}ڗ���1�Ϊ��S(�hG��;th�b�t��uy�r�|!-���^,�/k��v�}��@��ǭ��C}r�:��5���W�,�:��i1�6�U�@Dxf�&�!ݘ�ʯ8�ixQ5�bka&wz5Zi����t{�|��a������/@>�|�ݜ��p�yYK`ܗz9B�^��'��pv��t�0��ќ�5m}���@��x9]����_i�L,�n�p��sP7b�X�;-���4(��~,ݤa�R����ki����/�����>J#x�|h�*�)'U��1��ϡvϏ,W1n\=��LQK�է#�ak&n�Ҷ:å�ժY��䤃�韩F�%� �d����Iٓ���A���$���{@,A�>�	Io���:=�BY�*#s�<�]�� �z���M�G���dI�M��C�\޲�2�O�&�N�����<0��8�'	<x|8 �͵���ZSAٽ�zc�X9�&eFhS �tUh=��]���6y�,��ׄ�U�z�u�a�~S���"w��,�o3�_�6��V+��ݨ(;Sk���1%�]��;�"�5��7k��sJ�9!�
�����"�2
zS��dU ����V�h�O3[�6�@�j�֡�n����S*Ot�`�uT:�L��T	�9��:��{禟��9L��и���_Ƌ[On�_ۻq�Ӻn���W��ҫ:;�V�U��6^���Ա��^FR���4�yO 
@L6�K��g�Ò���;y@�m3E��j��d9�EƩa��>/k������S�r߄��n��Hm����n	Q�݉�!	��R)e�x�@O��>��4E=����jY9�;o@R���7�7��Ө��Y��6�/ǟ�`��?"�~ty�f�bV�	��hˢL�.� �?k�����<5��g!fD���%*�mj�W�Fz�����w�e|��bA�5(C�L^-Y�H����\\h�ڨ��(9Fߑ-+�f��m|he������OZL�y��M(�&�j甫���ch~N����C���\\$��\N����(*�uZT��FU�.�"��J?��pC<gT�h�%��W� �Ώ?9�u����p���JJ\���
`�ᐚ KS��^
�l�����1������kK��d���$D=�Zɐ";�H����c��y��F�D����k�+{f�YH1��{Q�����ÇL�����w�F?���#?�doǶ�.#�H^��֡ˉ(	�9ܗ�*�Tg%nkW4��N��:4t��,� D-$�2�K���R�uo�X��fo_<`�2[���I��C�Fg
�V>zA��i4�D���=�8��EjM������O.wk|�: xpU��<3�-���~jz�?���o��>j�@F'V���R6#L���ܓ+p�7��_��.�6_�d4�p��t�(L�o�!�����i`\mhtМa�v0h�}���Y_���=��El��D����Zgm�(�����!u槠N�?gI�{Hx��w� �@kB�;�U�yv�^�����}΂~���q�������"=&X�瀲3t����*]��΂3�G��������=�MZ�Ǉ��v�!B+�L�ma�ʔ��KZs~�	h��4��I��Љg����;���R������E3nnl��E_=% �f@l�@3I�G"���]����i>�8j�a	?���5Y���v�Xh�Gݙ���^q?�����F��>Of{�����Ds8��[_��}1T*sXP��A8P���C�Q���&6z����-8�=�Y�v�ǐ�h�#1m�C�����F�ҵ�o�i��@��C�Ց��j�5���7c�q���uy���0	/�9����d@i\��M���H��bY�Q>b|0��/�>GY�Ϟ�ʍ��[�N�o6ރH+K�HG�i��XZ+Y��>ݬɤ�n�Bz�� �܆J��%��������G/vJCx�G$�_���^}�� m-�֮-�0�Fv��8I,�	���A��p�8ȝ�#'�?_Ȍ�v�txb�QEI�K+mn!��8�/j��ˏ����uB�g��fV-��w��n�{�V
�֘�x�oO��C�,��|���w|�5����	�T�d^��㶓b�>��t��Sm��>)��&���f��N�Z���<�.�,�\�w�O�M����7����o� r�����R&���^�?�w�4y>��,����f�V�!����L����g�g�Kʁ�W�>Ⱦ�RI�zX��'���B����N7] ��K��K�A*�f<֦���4��B�4A��_z� ؟N��"˓#�U��(�&�K�ho���Ӯ='�w$w�)�*�ǘ�W��&�G�$,}q�e�N�*�'x~�1�x[.X9G_�On��oz�d�g7�E�0����@��E�Z�'���BC�:}7\���+{�f u�]�zi�r����C>�Y�6�����Ug�~J=N��Vb�5��/̿�W��=h�+Z���S��9܂$ ��X���P��t�)���d)��[W��(̙�Zp�g�O�?�!�r��u��m��OnV�h�]ְi�����B7U�^'�]y>�9��Sb+0�^��j��_��i��m���s���F$�~
H�{���X����R��:��$�������5 ����'�p��f�b:'�Ȫ�Pa�kp�v5��=A ��H
���+���v����I?B�B��g�r�ͯDI�u����AU�G��Gg{k�
�8�
^c_���oR�;ѭp'����8-���Y�]οx�x���!o�͐f�7�f"�eL�<�j��1���k	�����ϸ��[̱'�V�S�@�;�J��ٓ� �������ppކ8�sʹ!6�Z��w����s����S����u��ק�;�(ہ� J�[��i{�M��������6�Pi�N2i�W'�lL�E�1���<)�gX�pN��8���д?U ��Rg�:0��CEl,��L��	��W˿%DL�Q����J'�a*LoIg��%RY�׳�7��`9Y}�6&���g���t�v�b�AR��(]�++j ?�1���O�M��@�,Xz������`	M+���%�����K�}�m`��`ڳNK^�?�eSb�PG���yߴ�k~� `�G�Jn�#U$�|4�;O� <���4'���ޖJ5s�"|�,BЛ{�Ċ%4��+j��ӹti;c�9��F�
���k�wl����'|9��ߧcW�a$&�S�'(9k{a�l!@(�G�Q�d�3���k͉|�ޅ% 7�-ѣu�@�Ҷl��权
�2]����ވa�̬f��1�W8}��AgQ����.��Q�eM
4�j�8���طӑ\a�E�O��pjc5�%���Y�,����uA����)F�R=ϫ�U-H�*U���`[����&B�Us@(YjmN�zNne>�e0�m�{yZ;m�bg��l.p��o���{
������'���I�Ko��V0����\�+�~d�ew��y��߁�ɤL܅qJ�s��Ft�,��e�;�)�t�g���]6�yүE�R��Lf۶h� ��Gߑ�"^fl�AaZ3�,.�D��8���R�Qe��a�V�d^�#�Ԟ��1j�����Q�&��+Tí�6�)f���[���y�;Ԣ��d���7c�2$����
���BWU��n��	�Npj�c�p/��t+�9��UA����h}#~\��@n-[��+�e�7c�c��|��`w�[K���� �!�{���<���s ���3�T|B��1ۓ�ֈJ^�>t.�-[cԥ��>��U519�K�K� 6$�: ��s��0����a��nɬ������	F�S���1�+������ ռ=�M�7�9z�r<g���;f�!:�c4T#�P�=t��� ��XyX.-
������N��m�`�)�Ifܑ���d�A�" �aLj���5�4c�})8d�vg'�L���k�g%�W���Rǒ͓�Q7D�D�&��YL��٦i}-��[�cԒ�k����h?�)�+ܽF��2�,��S� ��H�$�YP�P��""�i�d�!�Y��H�s�`⸔�%��9RG��Ilɨ;��f"p�^�{�|��M�#aN�����t�����⠌�_�Q��Q�M|
2�{�_�N}�p�MS�<��f��.5l��`���A��#��FK�ţ�z��Oo���u�g�v���)K�
�pp碓�3����ҩ��)l��,d����T7�m)2�"� ��%��R�Q
�_&U3���`S!� �D�Q˵ڄ�ZS�/|{�e΅M� 䵃n��f�[�Z��D8��^N_�4:�B��ӣ�7-
�R���_�����A����+dX�3Z<�a����E`F�ܝ���e#a��_�y���5��8j�	�S��6΢��Hu� S4���J�'�,Eƛ��/�5�JuK�����b�g
ݪ��G��3����t��b�����e��ks���䘠"��W�-���E\ǻ�����b&z	DRED�t�[�FRv�^F�4��Z��C�_�o�y�oqR�Zk)E���a��Պ���[^.���9q�D��~	��&��!����f�]��F�7�ӭ�[�aф���E�3�P����,�t�s&�xT����s̠�N���$�^UEaxMxsvB�a�BV1Y��Wr��
���i	�o�[S�r1�`j��5��^�Ҝ�oR�MCJ�rh1���l��}'�`ls�g��M�N-��`�
���x3S�S,��n�y3+��.�%���C�)�����RP��O��	�[^+u�� M�P����yI��� �y5'>��ܙ�tG܏J���/+f�5~��;LZ�<��x�;���0m��Ds9��`�\m"�an�h�$��\�I��&!IS��O�f���F���V���ٴW����Z"O̹�O�G̋d���.���p�	8_�GH�-]H�����{�^����W���tQA�W�Q���J4�b�Ҭ�&�JX�w���.G:8� }l�Eo.�o!�a����}(����݈��'9u�4w�]b-so�Lf�1�"�y�Q�K�jE��y�xYH��]~��4��"uSO�L��LV;3��m�'�3īd�<����ͦA��\O�����i��c7�0�Ge6f�W��-�blt7�t6`B�'-�CP������T��������q�y� ����`��S�����LZ��R�9��2��#���� ����	M.��\;8�������a�V�1b�@S4��03�o�"��@S�o��(�w��ҿ(�X�bF`H����B&p��\�`�}f�W�]��钴�I�Pi����__gfMɖ��%�N[�.�7
�7�������ۣ ����<c��5F.��������I��z�M{L耊M��e�]��lX4�E�y��/Gj�x�J�Wǧ*�.�^`
ě�%k9�e�u�@^�}�ʘ1]>b�z����w�"g/���qAt��8d/��ϳ��d��qC��QR����zP6ۡ�"^�&��n|,$�HHp�=a�w��-�����#ƴV/O�e��
N/'��e��vx��_�)J���s����:�,�]acl��04�DI�VW�Q�)�f�6�|�.uT�Яj`����\����-��A������>�i���Йi�)(˨7�C�-���k*"JRi�J2��L&�5���o{�$���?�����8��Vk	���Y��V�W]6 7+��:�zt�W�~����j����ǈ�i ��S��ɔ���<�u*=5��LF�u.��+�����d3ٖt&��]A�r���t:Z쥟,ל�����Df��Z�[����] ��F�������#!�< E��Z���A�y�٨
�%��2v���/���w�'gNȦJ�VY��i;����ѓ��T/"W)�.��B~�"/*4�[�W���X����<(�dڏ�68E��t��+��ck��G��(5��u�3c]��?֢�wM.���i���J�݂�o��c�k�0�r5)u/u�_�薇���8$眛t;eSK�X��X� "s�o}�ջ�B_���wUd{g��&8\m\����w^1��Q�(��]�飳�w϶��R��������{蹐��,-����n� ����N02\ۑ�'{S�����9�;GF��3�SҞ7
�4Cj4��k�@����b�#ݣ>O�p�O�o�S��z���`�����rJ��*��z��b�)�aHr��_	'ܭ*/��9ˮ#�����˸��W�7~mc�1�k��WX��wO��©�N-(9�s���/��Y�Hфv�fWU����x��&�S�i��'��{���hT������Is�gf��I�)➤7^v6��Hn���jg�no/g�N�	��4gm�������PK�hCq�{�L��Ӽ4߮���jo��~��_�Q+n����f׮����k4MiDW^
$_u�����ہ��@/�*뜴]m�|ԄVe3�,	W� b�ӝ�����0�(�V.�� ��E����s���sZg��В&��>��"��r�"q�`�C�L��T����ؤx�
��c���Q�y6:N�,�_�K:�ns��Nn{ �W^㋀c$/�gѦ�-u	!�+,_4N[��4�H�ˍ�AG�Ʋ%�uPK��o���oG�w�j.>�f�f��8=v�34���GN:��+0�����'����U{���)�hb�(�F�9��_�)7_g;�Z0u
��)4f�11�.�����&��5��BhU�	v��9���!ۋY7%�6��ㅪ�����j^�C3�رh���m�#<��`ۙ�"8}w�ij�M`����%>��Yj7@8Ԭ����E����:�ͪ��`��3�җl�P�.�J����~4[���2A�����a�t���{E���������n;6���}�ro]�������I�_;%�%L��udP�k��0L�h7�s���ώ\��j����_�np7pw\�#X�l2�~|���H�� 2�)E$��"�,iڰ3C��2�L��{˟r�'���+���k�15�;�7/�K�Д�1����p���A�J�	�=�a��\Yc`g(��YH~�SF��/qD����)�lA��ބ�a�G�h�ޜ����!AI�Ȍ�8Q/}��uߌ�&�L{�t&��A�6���i�z>c�TTѾ���yYC�z�������,��T��F��E`�TjD�|������d��ӕQA<�F��<�e��p0Q��e8��8׋[@�\ػ|V���A����Q�G�S����;���H^g�K���#Z@!�O �#_�T��͏��LZșE�<�
�����^c*���IA��8�':l��S�V[���V	�vk���X"@��+_��sv9\��sfh��d-�]$ql�RL����W���S��ƁDavp[D!�r��>��j \��Q)�"�*̆{1U�hY�����p#����|jPf�]�/4�IQ�X�_��0V٭�1>Ps	{��,����^�	N�Q�RM���`r��A5_��"A?�I�me����y�r�}ۺ�g�"��>�q��^�Q��y�����p��]顉Y���&��2�[�h�'=+Q*�a�K��Iȴpf�Hi����Ɓ��������[�(qbD��@X|�}m���9nZ���/R	ui�����F��u(�O�$���:�xϐ��l�������}�R�d���]�d�&�_�L�x���Hr���e���/\5�����^3�CW�U-l�y�ȍ��g5* �0L�ɋ���]��f?� ?��j�]�s�A?T������G�o�Of�SF�l��ؘ�
����K�sKO
NF������
�l���3o��Q���L �MժҺ���`���P@0xi�Mh0)��i��K)��Y��f)�~Ȏ+�}��c��Ր�&����a�S�0_�\k�������e	1_E-/�W�ou4gԁh(�GX�VB��5�m��BH[�}n��Q>gE\�w���)���I�2��".$h_���3��$���;u�3�O�[��(�
S�ÕJ�"�j��iq}�]�Y�&,0��y���Nn#�AkG��Cy	N/w�C�Ѽ��qaN�'�$�ʢ��\O�8�Ƌ�%y�N�ߍ���먞d$x	��ϜhH��Um�Ov�?0f�}��&!A��"�3�Z�)uH�9��`��"�A`s2^S|����Ka���8��0����Q����El��r֙�_�e��d���L�{<!.]�B�VCl���xo��a�?�Ɗ�u�:zl�4|BQ�t��p�^X7![��O�3�O/�UA�aP��E+w����Y[g>�#�F��;��|�I5$���sq���s��&�V0T}F��B��H0l��B�1���mũ�`<s�`ڧEiΪ)��EP\&I�����ތ����n���d|f��؃o;l:��8b n�yh3�2��1���q��1RJ= ���T�h���c��0;��L����Z�V���������-�%�C_�*5��,7��4��:�:�2�Uʄ�פ��.{�b�V�ן�~jh��{=��#K9E�W��K��^�E���)�h?I�j�.(���h'T��V�v�d�H������L���Jb�iS�(_�\��^#���]�$8ߘ�B���aρ8HY���ޥ�7���%`j����J����zpM���9��f�bǏ@a6~z{�_X8��|X�Tݷ�Qm��m�vW�v��^�.zwh�����ޜ��h�� ��'Q�Gd�����~���Zv�{���6�'$�����?UN+�Zz�h�����?*����B}��q��N2C�%��[�f����.�XĘ�iA�e�o��m��N��
p�c
��ҍu��o>�G{�sI~q�i�=�aS�ﴪ�VWKеd�j	�d��B�T֏(�,��8�B�>G�E��j鷝/Z:D���ã��f�[ ����»�-۽|;��qѠAJ%�#(J)+mG�� �|.K*��9�=�"�����^�f��-�O�т�7Xac��o�Rz�V�I]R�M���{Q�`DxӚ��b�m!\U<��c�TN��̀��Ga[�}.�6�y��R|�P(k�����%g��r=���@��B�WU��q"�eR[���T�I��2Ԁ�@���i<u}4D�UZ�O
ӆ~h��4ll�r���>M��8�!<5�=������1��s�eF��v%q��)j��n�Ϊ���b��� ���9M��s�X�%������^'�9)�mV(!r�o^*6K��:$��K��;�������U\��JB�^}DYl�@�����^ؿF��vy���;Ėwz�M�F��B𾻯1	F'�O�qM�"�т��z���.� �y�%��R����k�ۘ��Y1�3��P�<��w5��*"L	��sA���A��\�LZ��HnBMB�ND�g��q���~�]e�dD�
