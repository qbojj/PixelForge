��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��Ί/���\�:��jN#k?��ʋͬMQYF�q��Q�F@���U&�4IZ�N�e�ʁ�hm'�����&is�W3>0/&�M�j^��^�|���+m�C�=ɖ����t��L��m����|gյ��+��ʹ�r����V���#S��V�]"!q�����Tז�ϸ'FtQ?�M�t���o��:X�9��tY;�y{5�.D1����{�PB�<��O,?\�"��P��=�\���﹍m2��U��B��#�^N��'��ή}Ÿe+��h! ؋�z~!�g��ӛ�s���d�	w��ng�ź��"Ȳ�:|Yk��o��Y)Tw-B$��uȇ�����慛`�<1]�n�wEus���vԊ1</Ԧ70%a�$����Qʗ�Z����\?:Tw٘��l�
N/܊��o&�8q�b�>��q�d�홵�����[t�ĥ���2�X����l�����햆�8���-W�LN�If�%����(�����_iX��1 ����*��:�Re-�@!��"��j�����˔=e��%-����Ñ�H�R#[�n2���������a
���R�S۷/k��P�B	��Vhm5�g���n�aca� q�$��l�s�����3T}mɍ���8/����&��^tJ�����-q[��a'ZV�+�^�M��}r,'S�����M���|N��n[O�]��;	�`����Y:����PPg���k	�����	M���֍���h.�W2&~m�	cK=v�?ϫ_xiU����ET'Mi�{#l	�{�|�C\��# g��cNz�*!e�ʻ}�Je�MzvlH>{�(��;i/�>������y`����?�'�H�� ��+V��vɖ�|wk�0=h�=l&���)���m���[� F�"z&7��@���8=6w�[�[�{�b��p��.�4��^����yy}f\ I�5�Ԝ2Clt�WA�KMA�|��3z��g#�5����w�o�j(��#�/���S�+�:y�7�p��"��St`H��v�,1[2��U{��*~�0���t�&�`:��%���-�O�^�ld�P��>�?����tۗ{<�	���53XC�.��?cy�Kb���*~���_ў=��^��K_�'�%�)'����z���	g�L�ˮ��㽔���K��ķ��I71�_�^�	�8	h�8�`�9�}#�Ŧѻ5�Z�"�V���mG�����Y�$\3��󺪺d/&��k�.�_�woR����B�ݪ*��6�(��Ѕ��fj%P.��y�zL	]E�����'J2'�S��Ә�I��t�����¢�q�񍡤�9���i�Y�[��[l�k&6ǟ���UNhr����P���,���"�d�b�
�˼_0��-�1Fc���΂>#��q���n�)��+Y>:����p`����fȤC�#�0O����*�#*����]v���<M�L����g��x	�[���ޛ��1�`ܻn�'��@ 7��H��lX��s�[����a�^�!����	 ����M�T�ݤ��G��<���^%�[��5�SU�ӻ�P3�o�Т$�#۔�Kg ���ݔ�3�o����zU��ծ�;,h@����n���^xt�_��'n!�[�|Ε֖�9�U��r'��YI�2<�g �u�MߩoIߘ�P�D�tBa�Y��M����D��M�<��R��F���#np�+\�A�}5�8�2���|z��Zx�.��/J�Y+I�"A�;�;�>����N�Sӕ�`�Za!c�SJre�1_��g�e��&��r~�m��jy7�v�+ >����ɡ�WuYl ;u��Cs��p�9]vִ֝�y��~��!0}�a�ؙZs="��}t�st�K��ʴ��%�<�K�K��3w��ief7��"��k(a�	�i=�I�@��3�#� �u~�ȵe�ך9�������_��:�5�gb�Er�)�ߗ�Н���m|a�Y�3)�Ҟ���hs�8V`I����x�K@,��2�ғ��:� Ｂ+6[>�z<t��<2����S��M��?�Y���\5�@>��$�+[��Z��a�=� ƚ �˦!{/c*	��I��"\ŔO�,�>�� �<�KF�q�``�ɔ��ں�[�A��~b�?8f���;�l-}fONX��r�ΉB����'�O��&����3�ѫ��]��ʺ\��L���Sru�Ǎ3�h��Y*�l���4��HJ ���o�i �o��y��dq3?��s�ƈ��L5����JA����\M���K��ܩʪ��x@]�f�@�����
痕�PJ���1Z�J��6��#��`��mM����3�씮#^��y����t�:�Ô_`�7y�4٘�8�z_�kj��l�:�bЀ-=��׳�cq����>TK�tx�a���:���?�B4�JG�P�{Y�hŦ�3�4>S�\RNj}
��+�.�װ��Ǫ��O�h��z�y��F���J��q�~~p�;����*�zB�*�!h��R6g/m������wk� Z�naq;`ۡ�O��qD�}%&1���W�}�a��U�)��H�R;L�����S����.��(<N��*	��l�#��-�,퉞�'��;�Rzs@%���z����D^�+�jҖ� ��(���Q�~h�+&�w�Y	��4߻}� ���6�}�,t��4�~�,��E���� &�f��\�j�K��Lօ�i�7`OS��̭	�!�zJ�!&��g�Z�."?9W噠M�wM'\$1G7ù6Rr+ޡ/h�V-ʶp�7��t9d=���
�����
�6h�_wB9+Mcf���p�4�@l�a)�,�Y��#��[�
�R�h��$�(e9��:~�GYt2%]n@G0c�#�\S����0V�M�TD�[r�n1��ɥ�QP�@����?dlyF�!y"Ϭ�r���ۄX֕SZ�_گ��S������փ���N�I�� ����~��ˈJ�#�B�;츾�f6ץ��M)4�������`Ei`��yr�2y�TG�� �֯*��:�'Wc��C����Z2��y�ZI�'��r(	r��0�#�bL8w��
���`�� �#�oeu������fv��.Є{�l>9�.^�	��L��4��U��A��e��G��y��Ry�sHݴg5��������-��G]X�P�`�۱J�А��	��������K��Rb;�[�G8���	V�}�M�ܪ9��M�m�e>a�6�=Gz��Ư~]�˺��s�ex�6��� ��Bwӌ�9w�[��pJ���Eه!� 4�1|a�:��yt$�r�T����6p����أ����d�{F4[��|�����d����t0b�s߲�>\��_�6J����,2}�b�!QHI��?�v�����Q!���z����\Co�4��jv�%��$�D�¼��Jw�uH�8������O��F1�t���,X�T��ͣ���?�1;��f����ߥ:��M]�D'������c.-�Y�k}�!G_�ަX��'�oo�̰�R����kww��0+ñB�P���?3��F`��B0?��ٽ�x�������&`>����	gby��m.N�&�긏�{�u�"��GG���_$�*=���w;�]y5T�~�ƪ�¯|�k ����Qn��И暣a����0�`���1�޾mҨ��hv��_�Y�[j!�Db��r�dr��g��^�>�?��(�`��G��r3H1�����|*ø]���������L(N~��������U�cv�V�huK��
�f��nv��v�{�^�����ʈ2W��I� U+h��	�
��팰����D���5����ۇ���,&6*������2�̮����%)���@a Ii�a'�Z�:v_�\��+�
y��:{�j������k��*Eh���6�2�}&-��W=�_�&N,�>Ȟ��&���� �.�x�8�am�3�]v���,�T`/�e� ,�/C���n��
~t�����4�?<ֆ�E�gz��0��>�QZ�E�$���<�A iȮ*��p����2F#�}���M��d�����7� �=;Σ�΄f�x�w���5�l�?�?NnE7�~�G��Cf�� t<�"KO�D��p�9���p����N�=,��Z#�}8�i��>F��c�=��f�����R7m$��`�������Z&�W�a~O�18n~�w�NS��\;yL�Z�.�;R�<���Ғ��p��5�4�DʣXZG�7�@�� O �MW��dHf��)����u&~�>_<�|�F�4�<���@�HD�N����_ ��G��)P���+��℠Ǡk8c7+�lɛ���g\�P��_t���l{d�3
T�_��^���h!�Ӗg��VTդ��B-�n@q�u��Է����z�$���Zo!x������1tJ���/���!��'�_�ۗx\ųԪdE$;��|/�LV^��� �]`^��k�؝��l�ʝg�3=W6�Z	�ih"��;�%)7z�N��HWDj	nL��2�����W���-����͍6Z���<d9��.�)��xdS��4�XA��_W��/�ȳr�[R˟C�V�O餭��uG�ך�+����?L�@{�k}m~�aa�Y���ko�>QS2�u��yi�K|�߼�@�{4�\�U+��S�[����V�uf�"W��j����q�ِf�8��������m�]z#����G�H��68Á��%���Qλ@%�`:�ma�XcQX�{#��,c��uC}9��c[���<CJ�%o�Qʺ�
�2��'C�Wٴs�Dx�+p�؃�Ku�s{0r+��1�&�xX3�����4$[S���U�HY�~�K⿢���ǽ�zEY��M׊�@+q5���^q�y�7�&!�A��Mf�������֖���tQ�T�`��O6��/�ԣ��f�)1��K��`� K��[�����M��s������k7��3�N��-?~JS�b��Y`�4��`�r��d�����Ҕ蛮���r��ts�0�ʫ'x��y.ٟ$?yS����8ۥ�9��ie�N�VW�]c>J����vx��N	 ��&�l� ���k��2��d*oY��(��:u5n��)�d���)fu�\�7@ч�!q��^�Q܊zf�eO�z�^���DN�.�)�س�9J���jqP���	<�+����SuPX�/\��qhm���n����m�
���XƷQ�yy�̹~2:-2��m#�D`�F{��+u��_^j-�^FTVf�h��:�&�+��%@��s0k>0u,+�Z�O�-=��_�l ��ba3���~�J\p=Io�#ӝo,u�M�ՅHO()�?M,�1��_>�G%>��tMUqυIm�ꏋ��R��!�K��l�e$5�Ea�v����:,M:�z�`im���}-V���D��&��&�r����j�c[�.��L=I^ӜɗaX��{�H4�d5M���8�6op������`&�"|zMNO���Y,��N����;E�ѣ>��W���@��2�]H��~W�[���l�hn�H�i���zG�������+�������ɢMy�I�Q$���u���m�ڑ����V���u��_�h�>����u8C�n�*3p�d�<o�'߀����U�Ȇ[V���~obP���G�$������h+��Wif9�U���L�2]lլ���dFmX��+�N�(&b}��m뷈V����*�?u�	���_3�
'*}_a}��d�c��(�D'U9�1^����r�sl��:xWl|,�EHvs�q���T岝��h"�����dģԶ}&yϣ��Y-#�?M����"�����kS`J��<�츘�;�S�)9��غlt��/Z�C,��j@�Q
��n�Sħ��׻��������NL��SX������}0��P�f{]V����nF��G�''/�M	W�#Yj.�a�V�/%�����4tAhT8~� xS�MҶ�#�G<��`]���~.	���JP�V�cR��f�>���ë����q����/����/ﺰ� '+nL�gz��*�M��s�ۍ�i��c�(d7������u���T6zJS��*��?�Sa�TԵo��Q�I�Cq�-e����e��z����{z]o"b,���Z�~�g���i�0��D1A�N���~��#���GL�5i���Ϙ�?� � �(����QYJodB_HL�Z(��η_&Y�l55����ޤ��N�;"S���������Z �㮮�h8���!Q����y����&[�uwg�ڭU2�d������u`���9w�̈́'/�P\u��;�G����l(��%��8e� q�u�x��-�U�ދ[��˘b�n�"*��"0g�No
�x�h fyz�i1��������	��(��y9���!γ`�hH�fZ��$Ҿ/ÈL�����)ޏG�� A7v����/���yrE�����Ԡ�u,��T.�x'l�N�����! �b��V�2&ߺ� &��,�u�}Q}�+y�}�	U�? �ngZ����,��6�	�a����Qؠ�gP�7�	���@�(�d�}���s��
*A���9�O��J�)iMu�ڌ.�
��_$���v`��ԂA�W.�W� ��߅�i+k���3�R���Xo��EV; �)�%B���0	�}�P��xdɵ���}߇HR	� �PI-�6f��h+��p�PL�jjmvt����g�v��%��Ǒ-���a�I��}��A�M��;�l��� ^�r�ф����gi�tp������.5$;��
]F����ˊĀ��bѬ0��V��)��xi��Tꜹ�A�8��J �SG���i�� �G��ӝLTc��8�G�=帿�އ0�0�@b�K�fC{F�,�6��&��4�Y��O�{�2r�>�P�:�B$�g]tY���O\UF��̠C����ժ�~��J ;¨ D�����wL�dM �i�5[�-Β��6VD�m}��^�`H��ϝ?M<����w��T��"��	�O�����ݧe>�ck$^ౕzW����>g��̡�g$ǧ��?�,k�����H���>K&|5S�"�t����-�\�& �#��p��-��! ,hjN�-���*�#�P��<	���P��^�i�፻Fi:t���#l�u���b(����>y�)�Vva�X�L�m��#�)��dP;�?�|�It�	�\@G���g�����>C�jB�Њ�ݔ.�K�6�5��|��-
����ńF�U��E��Om�6��TWh ���ѩ��B���>�@D�}b@�{� ��Ѯ���Mf,�e��� >n�<u*�?�Ă׆�di�oT����U
�K�M��O���F�=TY<�bH�m��T� � �I3m5����B�3^�Y��C/�qK�KN6�Z�FkVy�P�3�/���x��_#��% n4VEfg�����c�B⚀��pW?���0i��z��C	R�5E�W���=,�$n��o]���D�*�oE5�4j�^��x2G�xk�R�-�f�@͙�8~�W�Ȩ�4F��O��S�����̐ �y��f|�]���J��C	��C��f�x�Ӌ(P�`؎��7o�-	�Qc�4��"�},�B)H��0�eǕ� �}zA�FM���\��2kk��b�v�c�x-Z��w�/���{��'��Y���C$z��ܯ�_���LSJ�j'̀z��"��gt�O:���	��"n�o6iR�E��2�w:�x�t�k�&"y�:�4�m���]�y�d3�J�$�N�	L�P��� ��N���=&S�Q�/�ǳq�D�7ݾ�����Ÿ;j��/75��P�}�TYJ_�V����yV��g��n�g�<
M�m�\��f���3M)�� ܓT�)�y�y���Ӂ�˘�xon'�{��#���<
��#؅�Wɤ��.����d���o9�Ѫ�μ��/�3ʖ���g��9�� ��t�G��Co�p��w�ohG&�6�T�H �p��;�C�P`��P�4��	�;�&�uE�l.7K�w��V���8{	g��%�f@4���ȆPj ��R�K�����}�iZ�41נ��i��]Ifv_������}u�����|�_XR�Ec��X����&�W��A�ɺ��*�j��TE�
�Ĺ�1y"�=�� 4��r�Xӹ�E3�^'����}�����b<+�5�|-��w۰8�T^='�r\3^���E,���QN�m���ceIk�琴��Ei�A��ذީ�C�ϙ��Ff�����aN���p�<I���9���c�1f�}�4���M�FTE���A(�h��RԿb27��>4,�)Z�6Ii�27[��7<������C3Br!�H�R�	�iS>�=D<��<h:�u^JH��C�~��gc�	���y��^����(��ֿRެ
$�>9��?�7
�\�8��?��;������-mQ�L�tm ���Gs�xI�"��A��K�i�� .Y�c�T� Fm���6YX^Z`�cD�l^��Ό�Mic�����C�^�P'�S���q��2Ɵ.�ȷ� %�jQ�^ij�>�o)��s�1Iͨ�DC�矊CV�V9n+@y���^C�\��ev��_
���^t[�D���k�|������N�l��|`�V�4>�(�J\�aC�O�j�nR1��&�$�����7�'�Ay9�򍊠C<��������+������1a­."0C����i�~djm��My���������O\�쐼�G�w��&�$zY[�?���C(���M���y;p�}j���h�[ TdS'��I>rh�"҇��5xE��w�(��-��Y�*,a`���t���l�S<�v�>G� �٨5ۉ\e:���Y����a��PI��yU���ٻ�����Ī�Ez���825~��-)������r% 1��Ȩ�J5!�y�Lhp�Jb��i
(���ꖥ���i(�u~�ƣN��V%�hu��P5���:�I�!�?8xʠ��>� �m�1�S��^E��ʨ4�wb�DX���3���с��~2O��=�\�����Z'�	��o��ݴ�s��>�)'V��{V^+G��{*Kg�L�p�fȰ��Rf��:{�\(�i�$�r	�fq�ãBP���%�#�7I����mC�=�םBTbE�r�u��
�Ĩ�,�p_�B�j�n���i֖��zN�Q|�2���0#��z:�n�|��Gmi��)p�Q�S�>��L2L����𦕒�ok]O���Q&	�1��W��C�[���<�"���2�
�6j�0�X��.�ѲD^M	ɻZ�3��0��"��e!����&f#�z�~_�JW�!��U���� {霓�f�Zͨ��Iݛ%���hԁ�_���<�d��U��t�=n�hA.��
�� �����O��a풶?j����+��!�v~4��ʘ1q���a�.�.�����G��s�cW^^sq�Ϧӡ�iS���I��u{*z��� z$CG���8��MSn����D����*��|�O8�Zۢ�%��_�O�)©�&� u�Mo����0t�7���Ԡ�+�NB�}�����8�]�lYgx:����P瑆_��c
���!fz=���-��iz����kN�z�)�79��B3s�'��
��u�e�/7�>� �X��3��;X���}Z+��%5�h@����H�f�=��r(�6֣ax�*�����B�"�hh��0>[-|3$�^�&�k�d.Z�(��-=˫����1[V���EA���K���'�����ܺ>b?��9�W9:\���γ(.�u��E��yu��Eh��j�"`>���0{^��3���I���i̒�Ť,��y�qb߃ޟ%�׳t�mK%�V���ו��c=�-@���~*3[����ZE�h��B���-���hpk�G����[��N7���2���z���R����ǔ���Yh���1�k��	�:)fcc��bqV��~f��.=�{t:�^�>����r��;�!�ӃM�^�B7o������OO��L���~G��'��oq�]�������#Sn%�f��O`H�Dxvw;ʶ&��� ��qLs����vY#p������=�]���?*H�'n�/ꬂ>��%#�z�����ڝ��\�cB����C����dI�Z���'h��:�m_S�+�ҳ=��,MT�,�ǚP�o$l�˦g�$�`�6���t{YL&���o,9@Z<�����3��W�\ų�����Q�O{:W�-������l����ND�N2%���C����;�M����"?I!]��X\a��p%چ��&�z�nf�}t��j�@���7�E����K�G>>d�O�އ��e�(;�􌓳=��X�
������_傾^J9�2o�RԔ��H�\�������l�BYT�N�f�3n�����'(�ŧ�1�b�Mo���C`��6�=�k.�ݟ^r�%���e`a螳cX�����$�#�I��3%RE���9g�f��W~�5�7�7�=���\w�(C��PC�!�%(HD��%�܌��RhM:h� F�N�ز�PHW� p��>e4�q�,GvL7w����u�=����ؼ�m�K��)�3/q�΋v̂Ͷ�+7���]�!���"����WC�W6*�rQ�����g@d���$?��w�:�;hP�)�p�u����Ϝ	��t�Y	�|�?=���[��R!��l������Ǥڡ��)_�2�B�>��dr2\��!K]�#\h z�N	��Cؕ�=a*��]P-n�S	��`c>��ěN�bL4�"C�Z+	�A�D!�|�k�>�����i�6* ��?��$I�]r��;�)��O�bGb���~��!ltx�Q��~�%�6���	f�_�ڳ��|{qR���k.��~���%L�y4qM�/��(Y�p���P[_j�^�?16�ѯ��hKF����Z�]������OM?m�S���SR�!F������>�Pa�jiv'`�~FV��v�'�%@��
�:�՜qW[B�?+Q���ÌJ������!����d��.�� M]��U������x#�y��@˃ZА�q¯�P\l#�
�����,�����4�ZHO���g�+�;�������fcU2���	�;���M$mJ[��C;Lm>����)�4�Z��#�j���pVzԞQP�O���	:����y�mI �����.E�ˤ޾<���+��֒�D�5�^NC�46�ILpG�Ȥ��ჹxv������J���*Bdg$C�CoG�%����Q\�Q@���~�2�sq2Kzv�q@��3:=�랬ɖ��'�g5�����X�\���iN�_ǋys�j�P}�b\s"Š楠���y嘟�[��hkm���O�Y>�
���gQ0�3�����"S~���0�v��Z8�3���V��<d���rG�~�}�3��pO`1���^'#|:ℜ����>��a��fc�ӭ[PJ��ʥ�
t��6Ԋ��۝<�UH'T���tF��.tuz:�����*�)M���a�/�@V`��o�����S�s�_d��r�E�V�:�	X��i�i;7��){���K���z��/�\}����q��`L�'*'�Tɻ{�?��:��@���Y>�����9a��@KG�ȉ,��M�;�Q�R�8='��lW�[�y[�NIڊ �f�#���!�� �RQ2�{�vڐGϯ(,�ζ�{�n��(�l�Ɛ� T���Q=����Y�;�X�<.ϯ�`{�֣���͓.��
��
�G1�D ��mLǬ%:�Dm��"����
խɴ�6<ί�j�c�Y�f�Nk���d�k>��� =��&�-
Y��Q;{�H%�-o��x0'�i�P�슏�&)j�G/C�S��A **�
�U���/�����e�+�4>�2TOR��\�WF17�1ym�LY�X4M`*�lu��g:%�Ώ�gص�T�h\��&�DY�NR����ؽ:���O�G!�c]P��P}P;�Ć�����5JŊ)܏�Z��l��ue"V�u��ۤ�����n_$�8��ބ�i4�7�l�ѓ��s)���j������a��P�����qɜ4`��d�_�����U�7I��0��vj�"��=� ���S�1RD��Z��T���#9d��0�$%��kX���ܤ/�|5.p8��~�gQT��/�kev�� ��Oћ���
��O֊��V�qB����;[�����no�!y��w��2�V4��6�>Mf�Jۛ��s�*u\�y�W�L~X������O�=c�#�)z���dG�g��������7��������/26�n� �^U�X�[[��[�����kab@9"Ě竧�d@�Z"C`q�;:"pc�b�}ܞԌpZ�
b��_�2����HA��yK�$'I�B��2�M���n���o[��Y��C�
BC0�ջx�7m<5���)�*O���|������"Z݅�1�oH�'���G��¨��t�L'.Ig�_�SO%f��j���mB�����Ih�e��d�%>}�Z�����%��%o�X��{@�,��o�h5~��S@]�:e�shnS���e����
D��4�F������Z�mA�6�R�0���� ���J�_#'ڝ��V<ܭ�� ���)5��K��-ɵY�x:���UA��8�y�47p��/�d�RR:�Ů�<8��������VKz�ֈs�>`+��e�AF�Gf����P(���T���� ���¬�ƒ��Q��y�L�J\��G]�B�Ȝ�9F�"r�SK�C��"��f����0���� L���j����O��v+��0�hҔ�-!�t�N�{�+�O4-Vw{���k.< ��������c�*���gb��Xc8�팒>�S\/P�
���)K2[V d4(kj���
�3Ŕ�X�z�5=3.�O���F]I&}��9�WU�a����6���s3%G�w�ZK�g:+v4�ŧ�ԧ�t�5�Pݰ�C�_`��u��K�B��|��}�k6~˸qQ�=���Q�w��]z^�)6�e	o��s1������k�W.2�P�R�l1vM�f�|������|�I,�T��i���|ö����^�+0nIݐGH�,�=����.�������țp�fh�ynp�8 ��C&��`���{�un��}F���?DCp�4�R^/~7WIRJ�T[Zly���,�U#9��m{���^�N�o|n�v��p�/�v��7���ُ_cP�nP��g����j&��Uj�#��+2Z��AaUːQ�j�)��
�cR�>x10~f�
_|1��j��s] e�����LR�eۭ c8A)��/E�q��s�3m���|��W�j��f��sa�!9��=r@�{���*��5Z�f�k���׋���B�1"�J���[��P���D�k�Q�>.�_@UO
D�j펉�Aw����k�jE/�^�����A�n_�Q���Au�6{��k��8}�NvؿPL ��m3���]\�3�1����:t�� c��(܈n����_p|�:R�Ѯ�OD���f���������|���"S�O�
���i��K��.����8J�.{3��6)��8�1�ѵl{�8���y�?i�ҋ���*�PFyH��FN��=L(�e�픶�}�`�'NYVJ�z!z6Ջg����ᡷ�/W�mtj���t��d�ϱ�F�Bn/��p����TI_�1�D��Շ#��o�硲�Eta����T:x.��*���� ����x9*�]��{07�mڻq20 	G�|9�@]�ԧ����,ϥD�(�v�(�.QT4���bc<g� 9]���ͪ0��:2)����d.���X!���v��K�ŗae�o"��&�J��٭m�zl��ո���|y��"�_)��ڒ��*?�)�ޓ~�PwI0�NI��q�>�<���½�Ҹ	d.��qE� ���x�ã�1�i2�oz�!m���F�8?�Ķ�ݴ� Z��S��o�A/d6�$�k/>�6�aK�1U��o���x7Bp1ȴ�qU1����Qb.?;��F�2����v�s#��[~L���ϋ̤����3�piq[c�D�z������T�^�O��Q�G����Y3��.I	��F�C}���"u}ݙ���u+{B`Zm.X��2#�b/lV&/�v���.�V԰D�`��r�ζ�Kw���� 0�+�����T~]4TMi�2F���Ng����9^9�X^H`�{���'��� �ϡ.:
��Yi�ͪ�o��eXp�D�I��,��<�Ɲ�����u
�מVY�uC,:4j��VC�6��&��QR�ۇ�[�,1�V�������G<E�`	D��R�&	`�B����]��pud�mI��Ѷ�%pO&o����r��S�����	}e_� �>N2�k��G�������	�@(���c�?�yj���s5�dh� o��\��r������a��[PD���+W�T�����f�[^���d��Щ�����$"F��t�f-LV����BZ
c~xX=.�D��&���8��{�t��>Ԅ;u+��Zy^Gk� ���R�(�_aB���-f��Tԓ�Y�?�$��kq� ��--a����іa�`_^i�A@`em��PM3妛���a��S�k)���mr�z]'u����]w�|t���]ke��`�~�3�y�0�ŕ�E,�M|�BY�N ���p�j�d��V-q|����=`�5zq"!{8�.�y��=[�8�5``��7�2~�����v�e��B�eYh@XR;_\��0���]o�S�.����x(�oR&�n`Q�Ue���\h�Z�B����ĩ	��S]d����\:7����Eo�5Nx[��<�:�4�iEZ����C���Ģ��u�B�S]�������p�&ܐUC@�,�Nk7�6w��q2(:#9}r�Y��/N�f��#�*��9�-���-�i��a�/?�g@��_�Ӷ�0n4�A~F9�:D�����'��%�����	��/rϣ���Ws��,N�\,B��t�)����ٺp-�aBi�8{��esxh�Z��Ҁ'2J.��oQW���:F�+H�����m��"�t���ßǄӵ?}���{@�5��uG��t�B���6�*i�b�m������m2�)J���@�ֺ�����/�v�G�S�Τ���c��M=�� ��V��y�>P�௯��/lS�+�4WY�Bq�g܏�Mt��/�+����j}��L]��Cf茇��lt^?{tg���R" �^n��^�7S �Zt��&x�)򫥡�b��m)�P��W�:$����.O~l�I��r��d�Ĩk[x��͇�n�^�eF�b�}���1���潪���$U��<�Ij�*u$�����^K�Z���
u�-����P֠���B�؁�Z�ɄM.v�ְ3�i̮�tژ�lw��du��O��a�I��q�pDz���"��qy�?w���*f�3��W��A��� �����3�g��,�y�����\EUy��.��h���Ĝ�v���t�,��	Rr��G�E���E����G���Z,���z�X4��J�Y
FH�H��{>!����cv7��ļedqS��5�c�x	�JC���53�����v'm#:yD�7Ri�ݳ)�}O�*�~���0Z0�Ąl�خd��0hN�#��4'�C\'�kX��M�*�"��$r�PGU�����ox��=��z��C�w���@Nj�ά=\<��ɷm������pЙ���%�y	u�݁ֈ�3i � �,%/�^ܝ��Fy���|��ls �j��I�����l="����5(��?�;����v�1��	㮅��s�\Nk�,����b��DD?�v4�XL��.�*������S�d�!��@�sN���h��W��=;ɼ�s1��E���a"/DN� �:1���M�^�h�"�]�$a%4�V]Y���n8�A+%���kni��^���@J�ɾFv���(�ʤ������+{:�r��Bx�u�9�N{y�d�m�����e��$���tʟ�hT�+��t�;U������[�+*�X���뇩���)n�(]-�<�k����R��y��Ͽ�OGJ���0YB��P�ֱ��mj����b�[������^ä"):)_ ��HcE<�8~i����5�;�kf��+�@����R��J�8'��`ԃ��[��%�GWE��ſ����=�L)�iOFx�_������y�2��N�[�c�64�"�K
�?;p�D�]�%��̶(�b��WʟB.�>X~�ȟ��#�͂�v�� �q�<;[Rd�J��pfB�tS��0����4�9k�<���2L#��y}e9!�A䕢cj�&�o��>��F��
��ld�s �#�[H7�c0�9g`�K��j��{��7��>�#\>�%
