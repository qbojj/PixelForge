��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU����ax��ޮo��'��1�ϗ�
��FŚ���]���Q���li�8��XnR��yR�ß��R��
J�b>�8��1�d�K(��P�[�b����� 4:�����Y�|�!a�r��ѩ�`�ݤ3-����
�o��Ija��Q�P-Q�o���3�� �P���k��P`�R��P�G6k	��~�͇�W�j�8�+���y���I�=��`�G���l��7�[�(��'�ׅ�Ȱ!z��On\��j����A{TA�pR)2F
�^_��Vmh�V湬�3�?���b A~\��"�.ݗE���$�%��r]Vf���tY̆��-<�l�!#`}c0�xMu=ѳy���庮c�I i��b��J���_<�iB��pO>�t���?�x|]�T�!��!a]fq��@Q��"�D�M�������������E� }���,���"�**DR�W���Lq�[w�h����Х��L����'�X�0u��<�`m�V���d���w������y);Hi� ���1E�e��'ɋ���gCYk��;���!�pd�R�����t[���?�1x�~��M��T�XS�e�sφ�[e���q�g�e���r_� ə��c;�s��YQR�g�+�a.��S(�|'4��P���3y ��,X�?d>ڜ��ef{KeQ�$#8�Z�Պ�7P3r<���0FP��� B��k������� �"���s�QӞǶHZ�(˭�a������3�$>�@r���vH�\��A_���r�`��Yu��I�>TN�+��jU��2\!�9˚��[���0[W��X#M���C�w��*�'��Ij��o�?,�UZ(G�
W�:b��f�T�⋓���ç�8pe��p�`s+S�s��"�y���=��!�t)3H��HZ^V���M�����Ms>�W4O��c�G<�Ip��y0�8��Xϧ>�f���)iH��3A���"��MOMF;��y�ٔ����fd��t*����� ^�S�@b���qܾ6&��FK�*��Jи���l�3��V}~*9 ��-���u�p7�(�G�XF�@r5è~,`ՙ��Aq�\����>#|��Y	�pk�r�i���!9�?��GGH�1#ڀ3��b��ڀ'��m'�}Jʑ�|$�|L�&�f'��;�����V��I��z�"��"K���z*/�[�����2���>����67�y�Ԅ)i7�={`��^��j	��5CR�F�D�6����e�w���Ǚ���Q�:(���J5�~�gEL�Y1k�51�$��&�*� ��{u�j����|V�]p��M�+^�n�����7|�ڵ��+V����in2�s�gzs�S+�&�R�Gp�]�mo$�ei�SS��G��1f�I�z\�w'R˩f�=L�D"�07�1��������Cb��|�IP�\�2�ig	��?1 �@�ؽO��5�~�Af.���*�>���A�$���[�t�{?e��;��:}kK&�,�~�e�c7��d[����\�)E���S}�)c�9��O�.p�q�,�V�x��Gu�T���b�N����6ˌlG��m[_a G�Um�h��1qY=�UnʭV�X�����o(s��pဓ����p����&~1��u�k������^�~�}�Q[�V�`���a��}��'0^����9��,���1&�o���6qjЬx�5�������b�g����������"E-�f�x}��
}m�����B���2�P�Tyʡ�[4��r�/-g���]t���k=n���h�&�Z��Ы,8T-��`��YߎM���\�9��^�'�{�{�0��Y���X�]�X|��	 7��7Ip�d��-=�r�i"��>�,���",��7�iW߼o�W�Qea���E�r0>�j�)\�u�G�@<��$|�dt����S�&M��b9�~u��/�"�v����gy����C�����ed[#kEN��]\�<�fCV�#�ԛ`*jAPs\��.6LG��c������Y�U���D�Gk�=`�yp}�K�V�phS��o��io�d�^��I`�F���J���2iԃV�u�w�@�ʢ�`���53%G�ϼN�'~|�S&��І��0��-�þr��Re
Z{
bƈ�A6�C�����\"�w��تQ�q��Bk2�h���ߙ)���ܕk��9wx�����R�ah{�
�ςg�$a��P��k�L�n��)�zRQ���G��9m?e�lױ�)����}�h���#�ݍJ�Jf�]��+�K��0��~�|���Q�
f�Dv̓)�5�i�7�Ĉ�I���F��_G�h�W,�k�;h�$�I�LԆ���N�<�.��sӽB��������0���JN
�̔��Z{��!V���	ca�G;�q����$zE�	��nru�<�y���#�j��,��t�>�E^ɗ�,[H�k1%�+y���i� �a:�y���W��"�'����&��s�8��_*��b��q0p̲���aPwC�?�_�T�ih������i����e�[&���7�¬S~.M@@����\���	���R���Wпџ<h=�v�����kxf��ŵ|o���h|<���� �sϞ'�V��)H	�RG�̸?x�\"mN�/��7ZIQ��|~�hWV����ۥhm�Ci}��#�KMt�ܬ��@1��pTS�������U��O(��1��ʡ��T����ז&��Z���Q�*4=g5����4q>�j�S�*)@���͡���^��~���sQ������G3��l2㡩Ct��;�t�`�3�N�= �b�7��M�:<�a�.A��O]��7��Å5��ϓ�3R�Z���U{@iS�� ���n�s�y���=��Be��l1�^�|!�Z3��M����@4���
�D���G��~��%9��E�'�$��l�~�_��w����}��I�/�2�ֽ)ֿ��݄�I�Q�2C�-�����S����?�_|��V������6�}}��e�}w�x)	ͦ��.K��V��x2p\����ȋ�`�/݇�A�Q�C��s��d�:�/ͱ^�����u�إ�7�%�`ȯU�^�V�z>٬�և+��q�5㥜I,H	^�E�	�Sѯ�	�p;�3�3�L������D���90�g/��G�`��7��<϶%�1+�$/�6o+y�S�}�*�ѳ�`F#R��"!�1Sw������u�oz��9�}�W�jP��,�Ә�����"�f�0��vݗ<Fx�_��;������u�"��ޟ��#��zv���������^�6���G� �<�zk����uK�U�.�%�27 �����6~l�j��(����@ɋe����霓l��F:��r5�ﱡa"K��W��^�q!Ycv��b��e�g����	ۛ��w�"�Ի�D8ះ��$��O$�q%�J�eD��~��W��R�&5�ȼ��}����9y}�8(�Jt�҈�7���H�Òp-HT�)��'
������K��xZ�����	~�p��&�MU55��%{��(L�&z����'�!��g݁��]��Í����%?�L�냳"�H0�l^�\k�2�*���K3�QCT:ݑ�4���+7���h��jgxc�VN0k�V�.������Qm��r� �~޹�G�v�ƶs�
ܟ���x��������a��^����̿��_ 4!0�!5�V
����N���������YTjK'���^^���Y�Ȑ���j�����t-PL� �ևK��0B�QdmG;�oj�H���0�ry���.���H���t$6�9�a���=P�n��B.��h��ϤC��:�,/�m��eǗs��*�dO}�P֒�O:����?�.�x��x[�'K���M'C�P+>��/��٣N���v>����Ζ������G`��z�0CB�Z�6��)�;Ko��X|Y���#���d V:/Y�9(��U�u�N��+B�Z����)yH�_*�V�h�Ie����C	�&�HR�*�*���ƅ3�}dN5@��_ｭT��1��~����/�c����>������F�/�G�癶V¼p���B��:'�^�r;���*�5��bI��[��Zi�x�-	&��
�+�R�;�p��� ������Yg���J8*��ԁK�Y����Q�K����
vnw�+#�_LB�6#dkrHoԴ�P�`��u����]�XL�u@S�
"���U���$G
���tʇq����ap��&����ד��&�����Y�5�u|����;�vk��w��e��4F�;��Y����X���'��<@P�\9�]1���BX�I��bjΎ��f/���6��ZO/y��2�!h�tm�� �x�$i�a��T9ҍ8&��\�M{�M4m�H���=�?W�q���U�����c�����Mi�w�5sz���&c����� |X��V� ��{HsN-֫t:F:hx��X1>&o|Ҧ�e.���*�Z��{��+��u¡yg��`�܂G�ر{@#����]��6�_��?����3�Z��I��j=������L�j�qv�8�Zm�j~�(fuDMu���R�;A��M�Np6^bk#'�Qͩ���N�gNu� Z�18A��@����<)�� `�a.���)�%��l$Qd�}_�K�_�?�3�% �Y������b�dJ1�B�&hm�g��l�ؗ%�W�@d�GNţ:��1`(p�lk�X��&�(0�ۥ��y���ـ��������+�%η�e��r��>�.�h;�U�֌G��_N�H�Bg������!���(�X�tY��
�$7�w�^�6�fs�AT��43�WҼ����QJjѪ���e��X��TT����7�hZ���]F�~���z�e�(>����C��0$�G��賑��C�*ͦ�'"�˾S�֭��gZ2�c���B�[�.�ǚt|��V�����
*:"�M����wT�������t���\���"��9���o�*��[��Vb4F�2���It�������:�z=�/��Y;��
�l��0�����Txc�|br��k��+Ker�	me8���V"W�a��3�}�|qD7�&cL"�6	�y���ȊpT2�˗�Lz5q��Ӝ��̪���\1hB�&�&շ!C��7���'�:XZݚi-wݘ̥�0��؀�y](����9�BB�;v�Y�>��M~�<<�$�\���2Ώ��!~� .��X��%9P��30̞��o@~dBt""��Yn�B���Nɒ3�-���o�[��X�fC���#?ԕ<;M돈w�Ũ��ũe���U\?�%�o?�E˂��Βj)1�LdR�]{�F�T���
\��G�� _
-�ɼiʑ��O�fg�OT�L@�1�Up3"h.��JJ�ed�:��
*��=3&+�ǴV�p;~��)��
e�JV܍�0�5��!�oski����VA]���7�6��F)�4 ͕�s~�*��5��� �f�ڬ���r����e3Adl�(5���j�c<n����O������i���L������Q''�X ��#(ļX� �Ġr���P�0��h:���<�[K�in���_����2ʅ���װ�ՠ�孱��;"H�G�,%��ʙ~���u����lp���*��7�\���;�X����qB�_S2B`���4��ᝊ{�f\K���$�T�9 �"�����9�up�~��'�R�ӓ����2�Y��Cj}R�֙�Z�~)��7糢�_�j�=bL0�mP-*N�.�ro�,y]�b������O�OYL���R���㵮���|=�(I������XtTOu��Jxz�p���a����3��p�+����aB0�0)+ߜ� hx�k$w0L���l9��.���>ݓ��LX8Q6R�Ā"�9�z5��'�i!���TcԘ�����V�V��"�FpG��K��A �k> ���78���kio!�� �C"�sl��:�8�^�?�^���	m���f߾� �K$�� �E �ĭ����;Ny/[�S�1@��V)�˗�I�!�ۇ��MqAx]�������q't��2��&�g�,�C��e��9Ȩ��^�%����H��Ku���п�o���'A%�K�(��8;m?��K����4b[W�^�� -;vWu�;0S'9�����<����_Ġ6O�%�שlg1wtr�����E� uAYN��^������S�T�ɒ:�ܠ׃֏n�oT�.����7 Xd9�%�y��7��_z���)��p��#�$�a�[�k�ԗ�ĵ�0o5"@�3F��3�;��8Gâ��l�O�%�σB`@c�D��I�y���c�N��$��͈����3IJ"���\���.Y�aj����y����c���?��.5��s=ا�C~���XX��0ce��z@��m��Xl�o��
g'2�˵pu-�s�s�N��֤��@p�NI�Wq�	;6l����@|.�Ù�{	��A��qd�ƃ�b�v'� a��s��,y�� 〞=�P+�1���%��y��߫��g;FB�I�[`���@�����5v*��0yH�?*���F��bN2�Za.?�1��Dψ��۰\�T��
���~��-ν��Ϋ��B��YL��ݖ�J����Aֲ�n0'���?�?�}�EU�����>�-n�K=��m,i�E�ߒZ��Yx/N$�ю,��`B��{xAq���ºlvQ �拑����Y�AO�ǝ��]S$T$����x��.�z�)�h#]�����AK�@^�w��b$8q=���.��*���[NP����k��"H�_}f [�|�eÿ�.@��,�77�˙ׂ���ѺI�o������516�i�}M�Z�!{��eީ��Y�%PѦ�%�������Dv��M���!�<��Boe�d"�	B�
�|#thyD�:uEO</ʹ�ĭ�R�7߉��xI)��T��	P���}+P@_�8��}k���n���T^D�k�}���0zH<�ND���ؙG��R8�Wb^��ĕc[���A"v\I��Z�
���Ȩ*��cل�i��·�b,L�)�����w.U�kɦ�Qx���st�8k�]�ôk0���C�t�ֻ�t(�k������qdtj��@�.�/��������~��G#��oܜ�
0Ea}C�xV9�Y�<�����r
BR���o���Y`o�zAQW��Ps��nl:MR�׫��U�T8���y���ye����zN	�B����uIw��.���]i���d���zʝ��V����	Br�n/5��ǫ�o��K_���\e^r����!oI������p��2n_c/aR�3��YS0ȡ���x�7I�)�*�L����_'�,�aÒ�y�� |'I� ^�8���^����m�&jІ¦XJ��F�᧾�n�G�`qW��"7
�"=�B��f722~�dYrz�m�,>1��*�]�
?�!`�	Y��қ�>�'��;�	,6HFj��Oo��,Y}���a��Y�TgO�Lo��F}�;`ό�L��_b�%��۰Sp<�A�X�_�P��@���[`v��/_nM6q�>A֞���	�٪�����.�A�{ް����L��͒\~>.��rȃ�=��檕��J�J��JāRQ�'[ue�z�	�p����i��:��Qh�2e}��$g�ȸ�_��B����~�ߜ����u��m�,!o+�d�&}�3�M�<�ۍ�W��y!	���_.u7t˛����.^GT��(��1W�J��:��?���i�٦p�k@T�:/�'J�;jR6�.\ޱ}k�d�+�n=M��}�X������23ڊ�0@�V�J?�q���9�0_�_ސlemb���R�Mu�M�Q�b�����<�q�\;��.�"VxK�9/��Ы!�rŭr��`[iv�i�kDTv ����ʁ�����e��@$�|�M���7�8�0V��Z^�-�RfB\KΑ��,��nބ���i8�A}���')&��<X��
�B߲ɀx���h��Ш�����6�#����|EY#�4O ����6�2�1�FU���0�e�ID�@��QSo���ٽ�ɓ�)����izy7��Ih�;�Y��J^��P��*d��|9V��`(��*`O��)U0.���W;�Ok��I�v]1�S� o����ab�/Y���*�o�;��_v�e'P�S�r���2�<PO\�n�jF[�~@��O!V>��*�,48[�l�R3�'�]Pw4ڎ۪PT��nׁGg����<Hْ�h�֡h�	I��Բ̸?u%�2Ay���l��k��I�� %4<m<q��f�K�$д�{��UXd-�I^.+͠D{2�e��N)j?"I@x=�+�~9�����1S Ke�Y(Ys��Kذ��2{&)�Ds	m������g?r�ݹ�էs���`� w�Ϳ���Q��!�X�\�$�9���x��	���>��rhz�4<�_j_aϠd݆av5�1r12����Y>Ә����*��"^�fA%��7�����CG���@z��s%`�[�{�S���o3��ȪCH����N���p'�̼�̷�%M����i�kR��XG,�q�'�Gd��d Ӳ�?�!�d�<@e�h3��-���W�)�Ղ����kw���T���������]o���"��$�U���<(��f�a���
vݺNƲ�$�%����w��K=}���=��d�)AvJ�@���6���O������?)1U����4�����<o�L�b��Sp&�{�4�it�]��	o֐��93jNS�`�'��S��}㮛GQ�@����",xG�D�&5��2X5/���H��S����� eŦ���/ph���`V@�y8�p��C/� ��XH=�M��Hm�%3�໓A�qz�nWH�4U*�UO��u�U�.�V����'� ���A�U�� ,�܁�/ɏ��U5��ç����90�O"�x2=lPὗ����\m�H=73�3���n�+�=F� ��e>/|9������n���c��..�������He�ZZbx����h%�~-�`���H�a��K;4��o���b�fMɊ�9�[���K��r¿�Ōq�j���M�����Rr��dUw+ܷl4��X�ƾ�!��oV�n{
]�*����L����=����P�vl�O�'�@����x)�c����-�h&��o���U��?�n��xγ��Noۛ�O�4��&�����1L��n�Z�$�.�հ�y�^�\�_�ɊɹAv�����FԵ�n��1'V>$\�po6@:R�s�8/��<ڄ��GjгȢr�oΠ�CD����^*	y�g�?�Nꃰ��]u�1�4�s��GEզ}�T�=}�Y�:����d;ǣ��?��n�/��^�sr�~�� ;��?�a8�û/O����ǃ�({$Q߀��z�l�e�r��(C}h.#�Now=�B���&�*e���3G�*h.m��g(O3J�;�ܖ����h�C��,Z�&K�ϕ�+I�R4�J�̍p��F�S!��J�T+��@�g�����j��MK�r]o����<m�7*1iI>���
�u�C~���;⦴�%��d�|��EP�po�?ƘAـ�
a���2��#}��֭^
"�kZҦ�bLf��oBK�ʟӁK ��F%˾D��kU��X�_�Sz䔎�\\�����pk."h�����Ph ��GhygI�\&�
����@UIMkJ2r��F�YlLZV{O��<a%��Ǿ��_�1�� z�\n���tn��*�Ɂ�Izﭮ|}}�pX7������a��渤K�s��Q�&� *��b��sit��.~�>���%�7s�sx�� ��Z��>�2&-���z�,2=��l��F
P����ްƐ�N�I6x?�
y���|D?�����Ґ����7��nFr�� +9�+28�9�$X����޻�`��E�h]�Amix�y| +�/���.Ż���.c�k#��Jh6��|�*�\��S����|�c��}�͡����{Ӱ��KP�
8����,���������ꍶfS�������'f�Sφ����T�_�SEl�������%.{g���̢����x���`��S꟯�C$��P��������R)#$���~�~\QO������Ӊ%b*dpC����?��6#�̘����������?/h~����� x�!���ѼW#&�{�t�L"ϛ6�66)[�ɀGm?�H4m���Ʉ���m!b��M�"`΄��FPX$j�9m��a�ލ�`w��?{����*̵��l��Bx��Mw=i
 �1I7�o�����yS�t���g!�N��p��Z Э`B��V�TP��4������r~\���y��0T�U�?��)	��4
�l�����y��$���V�UA�����X������Ή�4�oVݒ;�S�GT����>.q1�,)�vI�pigi��;�<䈦�T2�e�#[�N�Ǆ�B�F(!��?$�u���D� E�^�m�&���{x����"��{d���8��FY���x�>�Y�۲�d���}6�n݆���z�{=X��"��Q�6�Ń~�LG�f5�97��kG40�޾�Ъ��ɯ��֩A{`sLyrE���:*[��["@p�R6Y�x��]�D����eF��@����̕A}h�Oꍥ�NzW;�m���^�a�I��j�C%
�+W�]�&���v�cH�D��2名j&-�[��K�1��2%�_�x����Sr�%�l"G���;�
V�=xX��>���
��yw�g�a�<���@T�Ҍ	�P����pf����H2I�[ ��cUu�s�.bz1ۄn\_�Ψ!s>���]��_�_U�=(O��<�v�%�?p�'�eY�T~�;.��R�����RfM�`��\ǙF`C�*GI��1�vM4�~hE,��T��M���0#	�2�b���써���|�i�-�����G �!Nq��)���J�� �P9w�ݥʹ�<���"d%q��*��w�S�s'h��� �P��ʉX5��1��hT�%C����mD,�'�Y�X�O���F�Q�8�]��U� <���{��[��#��,�+K�U��L�G�`<WY��rp�^���fVT��_ps&%f��y���5�D�:p�����zr,�ߊ�5�ژo0�@!1wx����}���R�7|�!u��b"��C� p��!����j)�;A,�ƴ���e���aǣ�;�b���j�APu����2է
��{��=@6Gw���~�R��	���YʕZ��PW����+��y����������Y�yr��Z��7�h+ᩝ&�yVKK����Q�����5�#�f���]=-N����b�:�_�x�i�O�[��1o1��r�-�l��>�@�,o�׷�0�?�]�N����v�c+g�ZC��Rԧ�	���[IB����S����'e�����87�C����&�f����6!K\�
�K8�� �8���u�i�ͯb�R�P�p*�*��O�|�<��Ip��-�/#�}^�m����?&�"�Y?�S�Ή�Yn�-�=��*:y���Ь�^t��{`T-��?���~�� ��EG�^YΦ��k��m�J���qU������F�^#�}A�}�W�X�7P�&�|�ڦ�)�Oǵ#�L�9�*4��=�+E2�?Ѳ�����<Tē���,B��8���dV�ak��b��4�,-ߏf�nc��H;L̥ p�t|=6�;1��΍���V��9�����d��|N1�5�W��Y�48��.
�Ԧf��	�G��OU�D��au��.��Y�x��� L�%�{�4������}�V&�Vc?�|� C{�5�[N!ry�iG��M����O��۔;t�\!&W���֡#9���F�>a^�&���F�����7��p>g*iy�;+�����$a*���i ���E�.��f�fX�V��cQp�3�Q���.;�is�W�l͈o��s8>��q?X�t&�������Dx���TΞ��hV�r0c����,�Y���tJ�N.�>x�N����
��$�z[��N U�O?�������I]d�q-R�r��
�V-*ޯ��-r�MB6Ŵ>������Ă��l�#V��!uHE`����HL��r�9�K{��A_�ӡS8���W�����m
ቈ��UyR���2�U<��3���&$�N�^R�,��Aa`�uR'�7Kڍ� j㾽'�k����>�U"�j�M/;���L�tK)���y)�������0|J�r�\f+0j�m�ǽ�O���������cq�(8����i9��HLr���3`喌i`ҿ�9�{�x�;���T���U�-�L��l�
��&>?k�"y���$�P$?���nE�F,��'��9n��J�9"kB�c�8��Z��*aO!>ݖg��F���E[|P=�}���z�����R:#����+��]�$_���Z����S�o��t�ZF� uBNv�bx��gLP�j��r�f15�Zc&S\����/s/u���-�H�v*�b��B5h�pbP���E�BS6t��DRh��	O~��l)ʝ��P��-�lϭQ�x��RpH�i�sD�]�r?r0���dN��MK�=�vn�\�L�F��T���m����Q;:����0eC-ij}�8{)����Z�u��>./3��;�H伩�D.��V��&��P�9FZ`C��� �!�ͪ��~�z>M\SǓ��u�C?��P��Y�qO���&S�[��5VEu͏����
qov�����^�m��۞AZ�|��z��/w�7fF�[F�5�x�G���õ��k#�h�㞲-_/:h�r��e�)�e]��aJ_ �Ϛ	Z�L�3uogr�n���Z�����e���=��ڸ�R;�]�g�K����T�ԉ�1΁�/���%�ϣg-�#PV���i�gJ����К�̗pk&�QH�[��yQT�Q[�~�fڗ;�\������q�2S��;�ݶ(��da4}�:2)\
���"�ّ�Ǭ_L��E����M~�n��';�m�*(�3���I �晏����2!��=��3<0l��W���R�s�I�P�D��:���&'��ѷ��N7�:���Ń�DH�����
��c�("v��@�WD�#�ݲ���"����n�kz�5l !օ���
�=l�`ֺ�V�O�f��$J��O�C�1N�w͏���Z�1B�KP�� O�����&�9$a�c�J{�+l#7��T��/P�AD@+�g���Ԙ=�^�����eŖ�)���E��c��N�R-|5`���Z��I��k�����1U�� �鼓
�%�N��
��bF�G"��(|(Ep�勵�K����J��긖��z��F�l�<����	�@M�	�.�]o��b�dһ��n�O�Z%�2�WbS��F����q+&`	��1��	��	��G�Y�B�g:����yL�P���p���>B�@pI����ؠ�8_��(9Hf��� q£~���bm��f(���-�+Q�� }�\���X�[^� �s5rMʲ_,����^â�d����ه�>�b��U-�*����m�8�"t/^�a�m�*n_��飘�N��V�qS�����2�n.�?�f2�!n$���� ���[���>3�X���fB�K*�Ǆd�PC�C|S!�t6ڱ��^� ���������k�p]�͖͟�i�X�v|���湻S�����_2�el6��3�f������+�u�� n��k��V�#a�(h���4���ޟF���F�γ��5s���5��X0b�e�\�&��Z3�����i�x�͒�R��
��o����:����ZM�A��@��>�F�{�Z֯��#��E��U��}���_��v�R�by�N����X�8 D�� e���O�9x�f�%V_�D�-�r=�0.�.�6d�L�4��^	Ga��Q2q���wO�h��oA����<�\���	����o�I���vnU-`dc��訶5�6��|�bSk�U��~��G�nhaC���B'.�B(Oly������������N����?�k�������d7<�EN	ߨ��
���-�~?X����W��ɝ����5�mJ)��N��Y���X3���kO�u���s�ak�Qտ>v&p���Z4��Q�h�Y�n�sAS�7���1�X������(j��V���d6n֠�`�X>��V��b���[���5���.!���GB�z���.dw 3��海����H�w  ��a��@y�;6ZW���ԕ�Ə.���o�4�]��B�аZIb0�����W��d+^]����NBM�D��t�;1�0+
�Ij���Q�(�A|J�с��C5V;�ܢ��o�)�ub�YH�{��g��I������<w�'E]��������8[�$��o#���
��_��HuNPS�ㄶH#�` i�5�b;����>t��g���� ^A���QFUB�/��=�����@�{�m�I�C��!������%���	C�C}1hIX�A��}���ڃ��8x���,M��Zy��ȰYR,p;��UۃW�����w1^���NW��K�=s\J�E&��	������!l��D��;�����@��.�0NE����d���w��'���^\E��ƈ^mR!�QQ�}IC�Wn�|?%�Q�.�HZ*1(~�٭O�y�I��d�Ȋ���6G��:�����Ӑ���_ޜ)Uwns�,ف��*�lN}�q���B���O�U7��G�J���R��8d"6�v����w^ r�}At�b�4r~��N㜡ʸ��C-�~����"V��ˆ����F�_.R�?�V��Y�����"쫌�O,��s�nl�d���ԉ(U� ��	��&)H=����ˎ\���).�SEJ�b�{[!w�P#���
pmF݄MYR:TK>�m��GT8$^ui���!��v��g�x���h������{B�|���K��äE{倩��(�f����:I�Xm�g�9��j..!�H7G�ƠMt�:�L�_{�O����y��Di��'���e�ɵi<kb�5o�#��̯5��F�B���n�
�>�~O��U��on�)x��)���էy�vP,�}8�(6m_����!�&4�(s��!��F��pz���"�/��Q� �ȱk$Hz�t�<I?��l�x\`9�r��hW��Z��%V�Ap-2EM���uG�K��^Q"�r��ֹ�9n�T�;� �~���а������� �8�J����*�\���f�ri����tN1>�<Č�e%�v�K;1x�������Z�@�-,����ߩ鸋�9o���m�Sn�G���=�.A#�H���y�,�D.���Gm���H�и�\ـ��bę��.�ܻa�k]Ⅾ�fnPQ�ގ���V�c��MC>U�=2M�DXn��M�ð#�.�|R�����9���ᩳ2��X�}�~艉��3��.;͸����w� �>�Mtk��;�T��Oh��p�-d7;��Ǩ��{��E(z#�gTZ�'�|�U�ch}���.�̐1�Ǌ��cq�������ĬSd�6��(h�f�@�֓/m}̵wl���8IX���&�Jee�}fŉ��BΆBhI�EK۱'ޛUj�!qa��D�I �<FU �ŕ�,��;y%�f�v��
Y��P7����P0����L�&��kO� �u�e�;3:�k�O�"��{XVGv�?l��.��)��x���D����k�?��z�km7�Ѹù����diH�� �t������F���^�Xy���"�ҺK������-��t�T98�(�K�PG��P�`�@ڊE�Q��R�jqan��6����gz��;�bO���_$���zD5\����:���8�~�2U(�����<$���EŌ���۩B��z���C3�+qc!��It�P_�_����كTu�<�/���~7���/���'Q�xt��\��j�2�
������:M��xk��Z!�>?9xO�x�G��r�b�h+
F��������e�]����A��'�s'�KS��T�j�-�A�8%g]�#�S�8���顂4��E�X��AA^��9�/Q({���,B����`,�&=T�L/QQM����܀�DD��o�xJj�Q��1e_�BU�6_Kt�#���G.5|
Y%n3q�bMZ���Y[���9�����6���A	�w���h�G�h�΅B?E�X!���m�M\ôE��tSN2�D�B�f���R�䜇��H����EI(�a��}��b��I�}�R�T>K�^�y�0����g"�_.Ѭ,��P6=t�V�XПDʯ)kg�>���3g�����f��?l���වK�*׃����N�nD��8��9��-����g&�!a���PV���<Yd��N?򲞲{UV�2���T5��Rn5
nZ�;<�Ү�_�9
N��'7ʋ���K��^��&Ш��u������J��D�Pׇ�&�.��Q�<	�^LK]!-�RG�?c6kA���v��i����Jvr�
��E�!��~HtҝП��T�r�l,�.^��c3Y�����~�ZXYc�!��s���Ȧ+w�� .�ߕëݬ�%0��h�A`���k�JCrcّ�#�PU��4���\�Yr��q��+�s�G��y��Cy�<�w����q��5�K�d	,��.ޠ|��vMN�1�}�c9�0BI�H���\Y6W�o��D`b�um��*T6��5Y3��A����ƨ�nJ���(��$�-�=o���� Ңz ��᠏�����:���d��h_�]9����M��U�k2����+!�r,G膬�� ��P��������!��+h���dBX;D0�4����y�ոơ�Ni�������%�v��~����<iז�	�x,Sա܍:/�7�&F�+���N���S)��gҦ��Z�f,������fb�&���W@-\%�Z`G���bp�x`;D�M-uU	\X�2�s�3}g�R�^��#9����s�BnM7qQ�Ԡ�
O6FM��P�Y���$��l�a��d��,e¢����&������խ�ǧ벤�$z�ɪ��Z������<pU�܀�L�g�<~��z�Ppm��U4��V��j�����+u9��Jr"<�vQ�w�d��)
���ܻ4�$��P$ev|_��n�P��׀���Q�{H���%�۲K�5����ӻ[F�YkqL��N�Ř�K(����Kȵ_l(>�h[7P2�<#Y�Q&d8%ܤ	^f��h�?X�bkE:����|6�ﭮ�j?�nPRB���_�C�0�\x�h��w8>
`&H}b���?����ݪ,�����t�#Jt�ڊ���bN(7�F?
S����KB�k.p������������S�}-�Hz+�Z[�<��6��BS.2�6V�|�ަYsI�T��(��v��T����@`�$��A?`�IATM����K�gU<O�4����0o��$���=�J��%�T-?v�I	�|���J�Aod�ZU(�*���e�?}<,`���νO�(���;�S�	O0a��H�>����ݯ� ����r���Z��zd��0k25Hpa�z�/$���p�@��L���e�m�qN�L��H@����Q1�0��/�`O5�R�<�EsF�B�haF�g�os���Ȳ"�p�N����8Ǎ���]]��ՙ�����]��FtU�\}Da��k���6 e�������ZU}[.�;�x��6��BM�]�"���ɎX\�J��}2��cA�ZN�Mق��&;P�഍�!�n��z!���䋅�q��u�Hfcy!A�ȿ#�w�%s�b��IX��B�=H���$����v���a����Ez�tz.J|�g���<�P\D�&�D��]H6����@{z��j׷��eg�g���1?tK����"EH�hFU3#���g�%٨_����t��*�	�UP�+75V1�e\������~���4���*RΘ���>�%$�v�a�>C7��\O2��P�ҵ��d�˨%�g���Cӑ�'%65D� D���%"�]��c~.UCXv�u��W;ċѲ��Շ��0"���I��Pv	�Yh��hGa*��5�1Tepb�d�h��G�=]��s� �P�XbN{�]7�M��)�Q�R@^�)��4vE�1��!u�k�"�O'��!�q����	�sX�)1���9�hn�ȏ��|���,�HΉ"�5d#f�Bq� ��?�{�_�Ɇ���qQ�6�/��%{��)�w�~8�m���
�~�����$^WL�J�������z 	�>��[�+�1*�D46U�n�K}őCэ}�������4T�3^^l=`~̩��5��.rP�{Y���}l�D�JW,=�ů����!/���w�.ǖ��;�GE�ӬjFgT�)��>�l��#O��i����c���4��(�8�E�l�P��B��TF^��9���b�{|]�Ԃ�1�*�� !���V)Yqh�K�a�ѠT�aۑ(��cve���h_���b�a��<����8�e�������̓o�@���5�/��pD�������P��ޅ<d��㗙�h�j�8[H�L,��,��l.��KYr1>���rK�\u0����L풉���4.{U��� -�R�3Vg%�9G���t���K��x�'
�)����&�C7�	 f�ȯ�k��j�z�6=X	��_#��w�=�
�s���bI���~!���֗�Ǡ^F=��xj��.�kM_ϓ>`���x���0)��͓O,۟���%��5�Y=h�z=�lO��9�#�Q��S�������I��&��q�Nk$1����{Xc�<k��ά��s��7U� DR����æ��hs �]��^ގ�@��x{���
��Lg$�N��M��]��$�,Τ9;\�L�_�UwᰢN%9+d�^�Ý�+=Rr^�W�)F.���|7�}3'ίQ}R�u�g3�ZZj��|����7�]n�~~q������@r#�Q�;�@���S����u��:��N���mБ��z�_D��F���S��(��b|�7M�༆�8�v�������DJB�2(�&��<w@��w^!v�+?�2�#����k|ߡ&ӡI��rk���2y$��O{�bm��y��0�r�ME�_�}�Ϳ.h�]���`�4LP�@0�_`���ij^C��JiR���^_�
�-M�n#�|N�k�~5��>�
D�k���"�7��#���p#�kY��``��`��c�wZ���$�
�ߨc�{��%�=�j(`x��EW�h�O��{����R9��!�y��h�ڎA�+��D�E�g*9�X�d　g��)�#9����YEf�����8�Z�o>���4GM������җyd�s}n�R����J�ܰ�%	P8iy�ڗ�`�>bd�.����@�k��2�n���EM�=�<��u&o�i�)�;�2��4%���#'ԕ�v>-p�r����sB���4��@�U���W���6Fh�N�A\�{<�5�U-�)B���"~�D�@���7�|�Ieܞ��,���}�>+ٜ'�:�AJ�o���������F��UTyӏ��  �]����eɺAVyȁo�x�;�{�v"W��G��?�����K��H�b�$N�NZa��aؑ�i�諆I0����06�ǞWr	y���L�?�|I1��
խ����U0o�b�R�Y�H�kUs1�h�y�3������ZmH&`%@%���(���#�E������e�\��g����5�ϸ���.�ƪռ��aƬtN�k��&A��S��)�ŠV6��M��G��	H�S�Wmz\?�����N���׮���� a#:TG�!X��&��D��k���VQ��s���w4rc��l<J8d�(,Zҍ�/,�FwʰG44/=/о����C'�3���iqڏ���(�6m��5�����w���jr���| �/��}�H^'�#�Q�j�����v��DeKi��HS~Xj�fӹ��S=/��=�ǼKØO�9���f���=y����Mp��3�٫:�ͯ,�G�^�҄R�o��[��v9o����-�7�c��(6�b�����+�:ّ���t~2�M�aL���/lo"�u9mn/fé�9�n�#��������v"��,]?K;{n��<����a�c��OFL��0�|S	���C?�c�Y
!ߞ�!Q��񁹃���+Dh��ʝc,/��@	���첣���G�AF4�S�OM��rxmE4�"�~7��~�Ŏ��z��$~Kp��f����:��F,���\�:���'�JA�|�N/S���f��Y����b�9o�S�!	݄�:╥�+����"Rm�R]v��V� �e�Hᆘ�XQ���w�4��5�zg%-)�j����N�5H �(8&�<spHt���ӞL���e��uab0�>3�z�]�
�io�"Z���qK[Qw?�����VѤ]hn*I�O-!�q
�Ʃg��I[�!�Z�������a��U�7��
����Z*w����z�S ��w��]�:Q���y��Z�����9��ֺ
�n����X�D�Lʛ_�.�t�3��^u�P��R(T�y�`��r;m�0ۿQl˓W�4$!�]/�hn3t wyt�J>�
f�5J�$��!wTX .[i�0q^�8u/��Ĩ6%$Pl��+s�vꝤe��%4��R��i���ŧ�$���0)Y�OS3���V��{>#�L�&>U� A�[���#ݕ��,M�o�] �@O�P�n�DF�g�R��y�O��^�'@��Rx��vs���!@QA;#>�Ze�y�Q��P���vR�J6�i�K��p8�X�Qƽ�\�\ڋ��[h��VB��?�����nj*��R 2@0S��J���ζK�##�k�l$��>UdM Q��)ֺ�,�S���K�_�CJ!]�(lQAa�ҏpE\~ ?�W�Q7�r� C
�w�������R��	HمZ�ĕ��j}=$H�g��?y
��s�oJ�>�����?/�tٺ� �P�i�*��8<7�A��QIAB��sR�@4+���h���Ѣ�x~�~��v!\�����
����9��l�7�V�>`V�I�|�-��[�ߡ"��l�e�( ���Y�Ti:e�9uAQ�8���gc"\|�N����0�Q��C^�x�Q�L4Q�K#�C��*�+�V���� E��Wr��Ӷ��k�?���7�tՆ�(MDk�!�!Gr;3[�������ͺ�o�_Ka�,�����b.VQ�y�f����6��1�j��V�AЦ여��x����X >f��AF-�⳻��2�"�?�1̰[���E��'G��x1�&Z��iv����ޛmם�d���]�������{�W��=��p}^og	�-�I(�5Qfb�����$�I&�BX|�E�w�c`���@��Z^��*����=�edC��[���;�[_p+�~��Pjm����`;���yh���s_Œ{}����Y����0��채����b��M���_�o�Uq3,q øJ)m��z���0�<΋ރ�m��r	av}�%�>p����r�Nj�%&ͩ��' �αw�FЫ޾���Q��$�L%��+H 21�� ;�ų}[��Sy�im� gP��9����C�j�EǕ���Mf;�}4�|۾ht�����P�l�4�!$�����jj[�9Q"�}�8�~�,�`T3w���h��� �ddx�f<-�JD� s3��.�W����|TEI9����KN����!��,om�1Z�#�*υ��@��=q�GV�uc�H�T[����m�Ⴡd޻Z�����N���"�d�C��T:s��Bܕsx7N�.p�5�����(9��:d�7���dΫ����Ԓ̃�s+j�#��9Ӌ��|�s��FG�V�=�ٴ� XM�%g뤂�[F��_en�vF1_�l�w)�-���<"G�k�4�k��p�����}©���Y<���+�J��b�=���OD�V��������t�&��XUK:�&dd��d�Co��H4���)M>��)�T�A�dM`�.{����Bm��s�>[�o�:@���Q�Mv߈���}t_#uڮ���#�[|Ζ��꧕����n�0�O��ҹy"
���B|4�_��p[�T;#7HR���i�⑲ep�tZ}ݢ�8�DV�/�B/�7�/p�[Qd��0����	�p\!��׋@f�1�|�±Ƃ�%��6I��"r�n���Q/�vu� �ʞ��d���^� �>:=m���O֨�/�)�}�I��������j�A���:"��4�}2���s�& ��Ơ�vfE���A���מ�9Xhǩ���I9\Y���j�ލh�1�V����<��ڜ��I_+�[lt`���U����Tg+z�N��N$]ʄ�Ͱpp��*���ҹ�#��r��P���G�#E�MzQ �<�9��u�̠Ͽ2y<�W�Į�۷J��rt��Hxܐ�#tp��]��O�V�5��ip���i��f���^c	��O�L���류�r��]?ژ\eŬ�3ԙh����=������((�s*F��\�I�?xͿw��#�w7�®���6>�n�,���}7P9��a��O��%��M��&���r���D��K��[YS���z�F�MY��8��� 3b�z ���}���JԀR��71�ы���4⦉�&��?͂E�H���uc�P�����|϶�t��[��Jǅx�0T^~>�h��+ǘ��j�3l��H�����}tlÿbY>��V���e�g�$�M�(���*|���\��Ee�&@������}Hct9Q��N��'����	p����z�D��W4�x��y9�۔FԞ��N��ю�L�M�T�db�}b�=m����^I
