��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��"�kj;5�9�5q/���"7ʲ�v��K?7���0�4�Wc5����[�ɸ*��F�SI�2v"GmC&�=��KU�g.7��-d�4�����v�O���j&��k�.��7x���
�n���F>�z���@�r�(��g�����Ȳ�`vĽ�d�i2���h�'��%RD~�:<Cs�fb��S	0PX�D���m�d��H��qO��ɾ�j�M%;�\Tzx*K��K(�aM8-\��)H�t�ҝYEWf�H�h�N�v���z�S�X�?��"�J���]�����;<�l�c=X�+���M�j���D�:��4�X���#)l6�΁u@˫ٺk���$F�Zf�����n����c��h�U9P͎��%#�]iP/�X�:����EI���
�x.�R������z}��)?S5=[�wv�|rҸ|U���TcHG�^�[�k_C
<��ش����qe�슘��m0�a_7οYR|��=�\uv<���[���]��J��w�;֜��D�%�~ħ���V�V5|��A����j�6�]�}�'�qCOB�~�\3���J�^�\Gǉ�m���PH;���ϥ�  Ƈ�`��g��W�;b���Z���|E0G] ��\7K�e~
���뼥43��Nt~��DJ���o�Vu�j���69[B�9P�I�k���FEP�Q��/���sD��Q7x��D��BX��Ip'͆i��h\��D��-q	7����|$h�Cp~ƤvY+U���I�#D$!5�'�ۗ�R0�� ��y�@�Q.������Y����wξ�{�j���7������C�$�MA���f8�%٫Sq�l�*��xO�����
|:bu�S���RR����K�*A�_��s�����R�G���$��XH�J�"�	���M��҅v��]-�z<���[ �N ��42�����*���RG2��o�Ǝ�t�&�͉�����hI"�ivVy(F��b�+0��kӊ?>}�9��
����u�3s���� ��/y��{zY�9#�/�8�jE���f���6�^��W;+��MW�2�_� ��[_N��k �Uo?�F}��e"����Ro�;�x.���;BO��U�s�WPiOz��~ݐ��j
^L	O��3.�juQ_��A���I)�]�ě�W��kjy�X���pf���z�9a��Cn��S W 丹�ǥ�F[JӋɖnp�u%�q��1$ψ�6f����p�o�O��T�e�����n0��Oy!�����߂��M�ƭ$�S�kET���b�("��_�?j�~��RX���^��|��9)�r�,��Ч�����`�-l��)3�"�!�U|���bK�������O��==͇�^	���ҩ)3�!�o�8l�5]#g'_��W}�#�Ķ
[�6���k�-�٫ꗗ���W��yi�M�,��'�ѷ'���V�$?&_�G�&=�wed�Ԗ=�Ҹ�"�s_/�ȃ}o�r��E쮤_�=^�RN�K����rce� ��:�36�iE4��֬���
���5�(P?���&�M~L̖U>�5�NXA�ڙ��ٙ|��~���D��I�B*Kuk6�=\����u�?��%�L����0��_�cf��3�!��p�z�5ƘݝP��@T�HDr�{��ө�Rp(��w��0�õgz�_�W�g�g�D}tF�'�):��OF�
��14�$�+�
�2L�z�c�Ǚ��>�y��?Ȋ�ܜ�o�Q�޸��~����(+2`��JB=��0ƊG�e�i����d�i�s�[�c@�D}����J�Ӭ1�zT�L��ڑw�q�B2�!�?P��ۑ\�&Z|s����y�I�0�ڽ�4?�u%uTZ�7+����LXIM��oC��9ꞧ3N�N��WV��`�q�u���щҒ�X
���%K�y����k��$�ʋazD5+��z@��0��߉�:�.m�#M=V�9�(�(�����+�5�5sf��
!'��N��f�V�4]���܎u,{��;��2���E�{/=��K2�ͻ^�<�a��Th(h�[F*�.(�ȥ��j���&��X+:����_���D��Ea���i��̲%�����ET&"ji�m�HI&�p�Hzo�OZ50��nӂ����h���\
2�R����Ј����Sz�3��^���;�d��x��<�)ё�Tl�,�K����MԿ��?-(/���I�w�}�#�����/3.Ӟ�B�X����@D. �s�^�#f�����uƋrI��$�0�� :+�
�#�3:��L֟U$�a�( �.]x}'ɿ؛`A7�ݞ%��Dv�t�٦��N�-�;�(`�^%iW����Eơ�M���xgJ*�Љ���W�5?�0ձZ�끱����{��(n��l`׀�G�q@K�'�
��R�zE��'B��9'�"�ȏ0����Fܒ!�z.s�nև��L�S�/��Y&_�
��j��t��m����.��*O�ޏ	���O�ws���?r4!�[To���R��%��G�(��%����*X�"O^k�}�6@�b;C5FҐ�3C3�-hb���7��-���E��Ӊ���S@\d���
x>�Vw�+�gd*�3�.���_��Sޘ�
^�(BG;ֵ�4_����խ꯶`հ�H�>�]� wg���J��<�Y����e�����=9E��KQ�R>y~���h���Sr�RNq'���i�;����[ɟl�{C�z Ʃ�Rb��mů� l�F����1{K,��Y�Y,8��(|�`����!���#�!�;�~��@��',����y6><�� �w�f���p�p��=l���"sPw���P���w���e�L!���Dbו�5�!堁�O���&'w���S��An���Ϛkcڰ�>��3#��R���D�j��B˞�>�-������:α�����|G�kT��F!��[���?ط��~�AiJ�5=�$GJ�����5�@��6	�t|����7�p?���oic�\�����);R-�\�� ��c��>��,~���o��sk=�T��h	����{����[Խ(���Lk�k�[V��\���V2_�Zy��#4O**��a��E���r�a8HZ�IEmR�|��X�A
�XU�t��o��.G���,��4����a��(q�����5�-W�JrC��[��e5��"΍��ܫ�	Q<�Qf���S�ۇhJ���	5��C�sm��ٲ���`!64gSG��~�x�0�����U��'jȡ]��򐣒�FF0ECO�"=�'�rq�.7������J�6�:�=�q�\*D�,�*�.���|H���`�x6���g������ƀb9�1��\&0�%���`n�x_$xye�N�(z�3����� ���:	���_f�lY�~7NU=K��Ģz>���KHo��]D���c�p�s��j�sXŲ�e5�`{��c�0H˰+��K�{l�����ELO�;V�LȌ�t�&��翛'd���_x��]X&��`�$�fQ��UgRaJ-2�o�ȯ�3�9K�'p�Kk�K"��� �j�
�Q���kv���;5d?ĎD9K��FO��������A�4�A�^^��	(���O�:㪖kZ������֏���#�����oW���T@�\�c�#U�����Y�)X�fР�:�:Ꚍ�̐	�;���8�H�
����P$iz($}�K{l %�v\�h�-w=i�Dz)U�Dy�]��x�a$M`.��eͮ3��[�R���tM�h$o��f6�1B�ҡ���8���խ�=���`4xo��=�H��Pٝ����=կ� �COc��k[���9�� �������f�w���#��0'������M:%d|XR�mCg-v�퓚fY�������\�l����A�ы���$g��Ίn$��)MY��m��K��th{�
���%2k	]��W��w1B�0EЖcÉ]2\��-����aH�)peU���'����4���k�sh�@٦�ߐ�VLT�H�{��������Y�ئ�_����<�I@s�?]���A���BI�|A�[�{ ө�w�&�<d���t׺}f����D�ƌe��v���H��&4�Vi���\�Yo�v�EH�׮£�S�c������T��}���R9�Gl֗��/L��5�P�j'����@��m�X0
� g���6Yl����+bi��!���rqH)�[霱���5?���3�"��2��-+ãr��]�MMK>+�����g2���C���{<�x��dl���0{�;k/K������\׎��U,�_5wDԸa��fF�S3��s3�1��<��6\�</�� ���x*��S�:�7�ݕ����T���@ݸ^	���yxH�{#2u��u��Sض�`�к{_b��:�E�O��zX]�����^�׹U����P|�jF�|�y�pQ�	[m3���{��x?��ar*.�ͩ�C�妤�Ɂ|���8W�#~�d÷ �?n�F�7��4k�k�T�Ϡ0�0�&��'���5�GY�U��'.�<6�"Sp��ܑ��a�[
?%J ��ti�c�mDɫa\�/�T��Wb�+�����NO�NM��ZJT\�Kp�׎���;�Ҍ��S{g�hK��v�K�[�EaAO�O��?�����k�Գ��e�x��BE�`�N�~@^l�+#���1T��n��I�1��.+B�e��bi@Yۀ`��bgC��pST�p��ilH�#��w9o�F7dz9"@<����5���q��>�=A���F�μ6�����,�*� ��S�M]�a� ��'
�IǺ �7A�lt�3�T�����tIȱ7�Ϯ+Y9�1�!��Q�`F��\����u��Q��]���q��흛^����ۂԋXꎚ�-�}�\�3��5\��I I̙,��t5��!M���>�D@{�k<�����?���3��w��:o�gZ�Ā	�jP9�9�o�YU��?%����SPdV����`�&�#�>���u��?��"	�î�\X�@Qh��&��~�nX���Dd�E�J4z{%�X^�¯��;���]��
��8ټ��K����I�)8|�	Σ\�'�R�%A�R��Q�Û]@�[8)�3�']�޶a�(ze�,|�Y�y� ���U͟�.g.* �rܡ�l��V����?�V4����0'�db]�xy�N��ls�UF�S�ϢU�! z����-�1�ظp��>�ޔ���(Cvp]ʩ{"��ν7ûm��Ƈ-��1/B��S|��h�OP�UNŀ���j��O��~�w#zxz��#Vj��y�)e��"�djĄ��+�X�A)�R)᠞x������g�O�VZp��FJ����g��2��� 7�/5�E~_�-�M�َ����]�*��(�����	�,?�[y�w��5��Z�x3���X��d�Yݎb���+�k�vlp�{�� ���;�v|� i�lAsAS�.�WT��V��ڣ,��D`J�?�z��9��*��z�V��	=2+�w�\�e���2�ɏ���Q�Xuh�/1�k��O����S��߻� �Z���x�X悍{|���4�C����q��2R���l@�Z3��{�W.��<}�lҨ\nDk�cJ��/���M���Ρ���	���ǅ�&���1]�}˅_N{�o� ,i���auq�c"-c���ۥ���&��׫��� ��{�w��4J�P�P�h��Ί�����)����f��2L���~֠���x�.������TM��O9(����%8ܕ� w�E�a!�P>,�� �{���i��?E�qO�*n�)�Ot�/Y.6(D+6f|,5o�d4e�<�ÁũJAau il��:6�������&�u�RvGhW��~fr�m�6�P�?���u ���'����U*���;��Y�,.!����˚������@����\���Oè���˻�q#��ƭ��a�$����'��^��²�ҙ��8��?ޡ�[<٬�=��Y,��O�P0��Ņ�������x4�={�������j/� Ag���Ce��Dn�RM�[�����J���� o����� ���VG���#6A����2��q6�~G.y>��=J;�k�R �Hm�t܇��6�U=����藥K��.&��/ �;Pop���N#ka-�Y�|ފ��n�0��-c��r��5	V4���(v�:�$��%�T���f���;cUȤS��iR�V@�f曲L.�A��fBCt.�$�"�fGĄxS��q֨D1�t5��Qp�����R�#	$��CX���(�6F��ϸ��-[�(�"�^�z��pq�~A���k�iV%�ZL)��ꄫ���"�=�|;U��uʒ�9��u�I�E��i^��y�5
�tۗ��jx�)c���&���6�/������s���T�b=�adK�U��
��p���b�|T?F!1��?Ӯɭa�+/���>Ωٕ
w�#i-6�fc�!M�1�U�y�;ߊ*T��� ��k!<~����bB�y�Շ�����k8��l^D0��A�?���W�)vF�u�A�;��ӎ _��/8����A"1���Q(�#�0��ǖ?�R���1�6I��ƑU���O{|�o�l�	���h��U��]�Q/jbDӆ$$J����.��m�����]Z<�s���D��ab
tt������Z�+�u8��&�iX-�/d�]�Λ���-���C&���Me�ǌn@ݻx�f�{-�1zv�I~�k���=� 4<��c��|���p��y�|_6�C�΃A��#Vv9�u"TfD GcP�����K�F����/S^	zP5J	����ƨ��ʷtD1�
N�ʐ��+��xY��ثi��G��6��� }���>I;R�ʥ]���ָ�U�����^��'���5��5wk��S�ϔ�^�H�W�N�q|���C�s}�|y	���wtw	0͞7پ����$��^{S��2{�5kϖ����-k� Ep{w-��ޜ��:�J���y?vҋG���<�a2TdJ�)ZgO9��ѨN�J��4o�0�=Y��ŎW�o+�y��Do�uc?�M��p��R�64�u������sG۩D����W�2E(�w���ļ�%h����&���)��s|x9�$~d`.�+iڳ:�����]�Ir�V�zyQ\���Su��#�PXv��=���[*$�������*�@v8��vԀ��i�*/W��[�~B�����kn���	h�� �.-��KV��~ZkT� bY�_Z�s�p��������=���B�v]ƽ���\�
z.���Sj���1�������:�y6g
x�� ���y��z�I:�v\�C��t�b���^كy�6�����2Kl�ӱ�2[�UWpE������5�
��FK,'VNu�ѱ1f@�|W�����n%?'K�b-L2Ė���ۖ۟�A:��EeOJ�.���΋��������	҄Kb��u�m�ab�/���r=b"��7zq��b��&]�g���6 (�f����w��s�n��_���q�~zcwK�ͤ���{n��"���6�惯�q�(0�p5�OY�)���o�#��q�����юO*Q "56�M@��zgN�p2����}�/����-����-��++
��p������U�|l��N�%��g���(���(1i��c�'�M�!���iq�����)b�jD�&�J����k6&(�+�e:" ;LO�-�& 5��gk�ǥ���:�]G�7)h�|�w��mlƑ#�䘡��q�`	���'������J��ަ��e��*�P$�1�b�0��v���a�F .��p���ֆ��{ń�l�'¾NI��r���n��O�jhY��QDW�����!��2s����A��>
�:��N�+I �e��P�t�"_ �nAn��*��oH�K�_P�	?��X�v�|�9gg0�w�@�۱T?�!~2��J���l��\Z"��9)Z�v8�-�1�%�����;�+r�{��B�+	ꞷv�ߖg�����!���z�`�x��5w�R t�mTO>��s������P���$;�n�b�iC��gN�j6�	ߺ�FS�����5Q�G{:�<j'8�(B}l�S���7u�]����G��c���\���8��E��4|��qU�zΔ�=�p�X|k�`@�Xj^� ��X�<����x�2o�����$�jo�c�Y"V T�Ī��0ℬ��_�	�%�)�X15�oUyE"��#,��4]�:���5��=����'�b�v����?�a�Zt�I����[��
��V_�Q��WX�ƨ�FO�	��I����al&
�/�H���TŶ���?�d��l(������d�\#\�@]�c?q�ŭP#�?;�ƅq�����^��yMٝV�����V<d+�+���_�d-t
�<c�_9>>K����Uk���nګ{#S���̙Ө�	L��7�z� �KL�x��'��j��7	2
 ����E�]#5��T��Ee��zuFe@�/v�: ����XI��u�s���Brm��RJ�y5W��AXW_OV�slAܡ�i:A~�o@��:8� 9\q`�\�/gy�����C���!���& �5��v��^��5ǟZ�U�,��7�I��o�$��^g�?vk��U�ڰR���ߺZ�_{�5P)������wt'd-���n-n��N�E��o�z�N� �!��e�Հ[�6��Ct"������\2��m�-���_ɺ# �魨���c�VJ{��{B1mQ�
����5�M1� E��D�8z��v-�ol-�v+z��=:�)����Y�^�Η0O�2�;>�LY?5��#,�I���p|��6��Z���!���o�lv +��v�ӥ��	�s��1A-���� X�WB�G��O:Y���~�g|��G����/�DF�@P�N����x<ai�Y��'�	�G��+�x"�	5av�20b��+�
/Jp�{����3?q\�c0a�hx�d����W�u]�E[�h��z������w�'�d;�J�a^_Wu�KzmH#=��)��ç���[NƯ/.�x�w\ps��_7,�43��+����m%���TG�¢1��4��G!�T�7Q�0;�"���ڧ�uS
~��Y�k��������h�?�b�k�s�g��������9��|�y�&�mp7�r��$l��e�Du�h��s�Nq�� 0fƴ�2W2y�B윀=���K3؃{���Xؕ��N�.7#����%��L��K-84ar�����]�|`����>G�zO�t���������gݓ�qp,���Z���j����}ZOyX���_�O���.���!S��8M I�z��>�K�`�#3���IG�d�}B����-��d0E��7;�q�1ڿO�ʦ̘�2��l~S���9_��zJ�72p���Q./�t]�Va�㹩�$���J?D�a��.)G�kޒ�_� (����*N�H˫��^#�Å�~��,>v71=��U�+ ��5
�En��(9$�+Ŵf�o�}&��ۭu�z�1���2��ȍe/q�G���1HLM���rM��i(�L	�'\�#����
2�����8�S�E�����κ�0��YF�JŦN��>]���B-���(iD=Ȣ�`a;���Ӓ���)۹ľ�(S�d��f�5m���P��g���Bj��x�U����Ⱥ�d�q9�(B�[����IPk$�{�s\�Ȏ1G��_�d
"e�D*h�<Y� l�0P����8�S��{�m���K!�6�W¨
�~S�z�K��B̮��X4����\��+�z��n�t|�f{b[ ��a��e}mT�W�.���/���&2��I�bB6�a����3���ۋ��DQG�O����k+DL���<�u)���czsZ��z�{�z[�8�Ed��o�p��t���|�Y`�������?z�BU��n��!x�I1i~����)�u��"-���*~����ﴠR���Z������9J���m�tE~<:ۅs4��7&��IO�l���&�ӛ�	ina�q��M/t>{��fr�e]!��W�W.C�� �^#G��Aʴ�X(B�5Rs]�!"&��XW�[� @r`l�D��D�yK���W�P����qv}�������6擋6S�*1�b�S���y,���w�+���8���T����f�֊`SƜ�蹲��3�]������nL��s~��X�h�3�'��=^�.�fH�d�� ��X>t=��i���y���ӽ����S+�r�c��`��#����k'	�!0m�����<�0��,8Iwo����?�bUxE}{������
w<O_�VB���ѓ�V-"��!�N�]�V.��?y��RGR��wM���N:z���|�({�U -_��V���:]�ط�]�}mǰ�2G@,q���D�++�Q�2�� ����m� ��W�7/C"^ތM��^�.;�6b����k��4�e�a&)���E�gb�w!faF�;ఐ6'��C),�Bن���1������z��)"���c�ͬ�W�[����j$@�R0Y�Od��7`O��/
���	�|��v��6��ָ�w��jvF� AIʯȿQ�q���	����,��L��K%4���2����=����/	��Ȇ���\k#��n���@e]��8��4t�H�&�+!_���=Cȩ�s�U�tz43�=��z^ѧ�{t�o��H,��`��r,����@<ZIi�X3!4�k�]@��_�"�
�)K<�)"�F��1�5}�K&�nd(�g�*`��7�Ɩ�q��іg�i��5�������Dn�w�<~��B�5������U®�N��۴e�D�o��V.5E��a�!UV@ޮ�v���P��ڪ�~���xA]A�U�/WӨ�&�łT���9+Hpgh�M�DqH�* S=�k_TBDn6%i�Z��K
��	<ܡU8���&�S̹%�s�(�~��Ti3a�B@��&ɚ���.l�)�����V��NI���
?$��\K���(+X7s�l_|B���:�!�8�(;$���-7=���T�����xOz}9D�9���	��Qrȃ��#J������^A�~p��܅ .�l����F~�p�"��Ld�В����	Z�\���)�9C�HƄ��2����������
�$p�l�<-e�)�fK�879�o�G�C��r꼾��x>B|Ќ۬2�z�΍�S��Y�`�[m���KCa�g��6��֚��\�di��c5� �T�z|y���F��u!��z���4�?�2�k>S�=�[�ƩF��.#$*�3���d��M]�	b���ɑGf�������J~%��s��@�<Q�s���=V��&f
:a��8��O�m�_Iz��En��\�DaMɅ�vHHie��C_�ҷ����,$�.U����&T���с�:? ����?m��@/�8Qpv����e�|9��[���8����%j�O�~�b%�
0�8�u�B/��r��4��x�h�j(v��U������7ڭ�Zb@�6]����:=���d=ڢ��@�:(�'���q� ��٘�o�R�b��H�����W+����t�:�,OGBZ�cN/���X<!*���C���9��HH�`fc�(�;ks�"N8�[���u���E���&F����N��� ��ɉo�㥑V�_;�<�>�u3�i�x&l�ֈ�-�	b���m�U��t�N�����ȼ8�_µ��O@e;As�6���J�t媟�m��&�������Ͳ�딣%e�	e�5���a�2�5e���&���H�'�ҟ�_�@$��u<b�蜘�L���cr�a�+�����a�Ǎ �$���v(b��v�U»ߋ/�?[f/�0˄Un'��K!*О�dӖF��0���XD=��t�>j	�쵭xG}��I���wdf�+[>��Q�q�6{�P:�ь~ ���O)�g���$T(���V��]��)��|yE� �K���+�d�3B�`��ں��-f>~�L��:e���dGHG~a<'O�bݙ��k�E<��<%r��!��C�k���גΛd��F��Ut�2�姓a2Y�=��E���Va"s\�
�tr���M���ӵ�X	`�xW�8���< 1]��М�9�ء71�G-a���`L����R-��a��N���������9Ih��fŠDN]�������"��G�c����Ҋ݈����Nd=LT���#i�\�rGpi]�1Չ�{����W p��#w�?�X��}&,l�Δc��n@nh��m�8�Z�3ʋZT��OC9�J]\J�r��a���p��/ގ{�!�c��s��\��?�ܭ��I~9lF�Tyޮ�΀����+����xSP�}�����x�<�7䌶2��ޞ�UMõ����d�����6��	�L89Y��!�������Z�� �c�3�=��I}���_	�����]�TG�6�ȥ�Q	p~��<!��U��;��$ɮ�Jū��}'͂Yv�vB��t"S�������}@�=���Z�t
�8.[�H�p�_�?�.kh�$��<�N�Ga�~:��'OX��w ~����j��4��S�O%ۣ�{/�8���uqD|*�X��DEi�"�����*yW瓓�X<���!SP��B�!㾴Ũd�f�S~M����e��C��A����������czt6]��jlZQD�zD���Ou��2&&��B1��"�M�Z+��{��U�h���H��^v)���ڎwv�6_���6�dq�ӑ��2�Ⱦ�ҋ=�W�tb,�3����n�[ޘ�xfG�7��i�sZ���;�@=G>ݸS.V旦N2�V��uBP̾�V�������}W�!��F�Q}�q�OP�ߟqHm��-������詤���,__�5�(���m��Dnp��⚬l�[��r�t�t˞���n&`��A���P}�/2�0�s��#t����Y_3�R�傝p�z�)>��k� (�7VA���fWrPKĭj[)�1�kJ.�Ֆ�#��Q�㇀�7�q����aZ����N;�m��������L 	�$&*#,;f9P'�Ϩ��6������Ñ��A��J�dI�Y%�]�_:���?���.��`�x�ދ�׶;�;�{������?�C�gB
w֖���Jf /<>�J	�o�Q2�=oo��68.�Y�ȳm�9�"�<��Cʽ�M���xM|Gɷ�G��LHj�D�j�.�Ա�����&��.e:cg�ۼ��ln7'����DL?�؊�_��[Y�(�e��+���m�m�gql ~��A4�Ǔm,I��\�hT h
�-�l&c>-3[�/@�rZ@jh��ryWI˘}��.����Y�#ؿ�7��P��r.(���{��<Y�����W(��`�����b8�Σ�p�~m����������̐Qg��� 3�����A&�T�V2/܋_%���l!��L�H3��2���,�C4�g��J�O�\�6O;1E��T,�wR��2&���p������U������+���D؊;�q�4�ӹ�`��r(��`Fzq�"���'5�מ�?F�I�ǎ����y֦<E�姮��́4a�#�Pi:�뷆6�0ԛPx�\]���2��������L'�>�M�Xy;�>�}�ޏ�?�}�D1�	� ��pp��#�xj\x���x��ܸ��sZX_{jps���N��:z^G��_*�jQ��TÉ�m�G�{��F��ξ�>�pg&�������H��v[6�ý!"BCNᲚ�_T������,��ls�#)���~Q�G>��lYW�'�{9���X�����"�	,G'�1�%�+��3�Xs�~�-�Q��r}��󸯦�� ���+P5T�'l��Yh J��?�b���q�껿�1����V�l��M�p���M���5��"S*2<"o:b���[UP>~*��(��+/��[�,�B��$Jݾ�t�����_`Q �[ʨY��
z�2�{1��V� �1(�$�;ɩ��7%�n�?�'��T������U�?O���,�:V�:g�"3P�� #u�xA�����#�aP`7��������h��0�Y>u/6�c/����h�یR�URյ�p��yLBM2�6kQ\"��qX�KbL0*:d��:9�^.���3�ّ�!n�}޽81-1������hi���󵯧�	�Ù?< �wN���#u�HwE}�"0Ľ�+�������'�f����B���B�Ҙ�Be��<gb(�Q�KL�L{g����+1G�� �@s��y��(��mc��d�Ǽڼ{%�z$���ү��g-�p _D�K�j˸��?�}���~47�����b��~�e�dA�HH�JRʂ�K��OK�o*3�>X�d)��U�� @�6�y7�a��Q��w�b��v�� �\ieOnY� ������Aq~�\M�v �`V���4o3&���rn7��������&����0+m=l��=��ԃ�
~8B���~Zn��ˍ���)W��xgj����;DSU3�ׅ�*�w�u�ݏ+;L��/�n��g�iЉߨ���Oõ����49$]gx˷N|��� ��E�RXK}���G�i#֨wz��F��|A=mcy1L���5�K�7��;"�w����-,m�ko�6vm1\=Ѥ�������R�Ƌ�985��e�����'�a<5��Al�iH�[D�������e�5�$�S�f�����/�`W�Fd���4s�ݩJ��i�#Zl��q���[�;��j��dX>��a�[�)�-]֬IV~/�� �fr���;��j5���e�	� 󌞘��wE�X󏩊��c��!�O�����p�ݒ������Ԉ*�]P����	E* {�;u���5sJ��]�hl�
"bM��jFeCǣ825�-F��54*:Pu28A[�����e���V7�y*nt{����f����'jnmc�R���=i�L�-�L��-���x[�J��VT�O�t��>z��_�ߪ��s��ɝ����O b�����*nk���%���e�,�pR�x�o�C N��Y*�(L��o0��Gn1���0�z7�w[���6�
�4u���f��ϠebvXaKB��{%wn�Jn���k!*at�
��,G������(�,2{�QJ����03�T=�fT�����Gu��>˛x\�� D����F�r��6�"�6�v��T�t��0��a�o�ZP�ZqVVF���G�G>�.�A�̄Xގ,�vꨦ�i�@�S���#�)���> >#�@`z-j�Aj��3�� `W/�@���Bz�̋
���ϺrE3��@H�н皻����:
��ƾ3�;�'����vN�؆���E8@ �U���Yq�V�á��܌��С�z��}�5m� 7Q��������H]�� �<�u��&�ʵ�Scrue�ZNkC2�rV����,=	z��$��d�'��v�U1���"�i5:]
A��PPN��H��u��X���,�g̹4��-�U;����^ ��}��i��SIx��i��n�)��w8�1����-�XI�y�^�㰿��`!���Bjfp��ߟKI���g�^�A��D������9�0\g�L�v����p���ʹ����T$�ѣ�i�Y�����!�Cg��u 75���a=��h��J�ޝGҨ�	�����C��q�e�Z�X��)��}g�4�i_�h.���Sv6���8����)�s���
p"�88������	Ǝ (\>��3�9�c�������5�D���í7)���c�r}Z��,��}
���C�Yڮe�Q�P{*����!l�l�WR���8�N/a/̟���zu��I����vb��Ĺ�F������>26�B� QӇ��ڵ_v�'y��������YZ�"�rcچe��4���F3�k���N<>I{b
c���ڲ�.)0���}�TZ��3�ҁE�*��� �3F~� �z��Bjuo��@p �~�YE���*�C��;��bV�ai�ˡ�r�-��~to�wX���9v����~�Z'�a� �h>Q[Z��k�D�� ?%����ނ*�
������˯dqN>B���H$�1o�y��4 Q˵c��u����}�F�@���)\�����Oܡ�:U)r�z)��U^�<��p�{p�zL�vx�O��@H�+S����P���X� -�Ғ��l���x�c����50e^U��28]�����?܊(��0�f�� ՚8�L�vCm����"t|Z��eA�$�P<Ʉ�E�T8%��泥�IK�)"���ׂ�S�}Dh��(0%�1����_��Cf̨���ĨT�r�(}ĥ����7�������$+�w\/��nh�BI�f[]�`hbj��jϭߜZ������󘕄Q����S�'=դ*�y�ﹱ9���4���{7���W���c4��9�xYm����^�Oe�n�S<�Y��=��v����,%|VPT�0Tѩ��v:9�����?����bR&�AѦ��u>���g��:I�$�
�j�&�V�p���r�r���V�)kM��Q�����:\�'ݺl�氋�,4�LĞ	�#Y'On}W�uzY��:f�ވQ�M�d˪��=���H ��2��2M}��̔:�E���w��Ѹ�k�����s��Șc�&Lӱߗ�ˮ����)�{��i!�S�9�f��[�Y�����2lQH�o�G�b<�qU�>�}���m�&Ц��}0���gz�X��A��p����{��O~���K>�ׁ$�	Y:���̫�|pY\�8.�%� ��at�:�f���+At�s�&R?����6��#�f,Hج���t�� 2�}���P�n�`H
���=��ݮI���l�R=TXe�������U��I�
<>7��a�'d���C�����"�c)�^؎���gѪ��������j��U6S�3`��C%���[b4��u��z{�pB�65�i��B"H����(Cw.�Z�׬�G�j^�sMw���tGv�M�W��Ⱥ��{��ЏyK��H;�tքk^���T���$�y�)ӥo�����/O�JD:�Z�����(Gj\�`��T���� }TL���ֵ��Vi��u:�xMS�1z�û��W8o�� � l|�/�Gn�
�;J����/�u���r�_>��~7�R������B	'eU�;��ƞ���6�n���f[��CV*��L��+���AYr�H��N�)�u� �eDq9���Д��q"<bxCJ��C��GW.� �r��\R���5���Hc���m4��T=h0{�O�5�����艡;/>O�-H�ATne�}��2�Z�6�+�� �x5e�#��5�FYB���2"��eϧiU.1��>�� ���e�S�����F�]���"����cjm�m�0�]Pe�Dʚ���t�~biR�4��̩j�t�SG��y�ˡR2��� b��ujf�L��fh8FR��?�w�$��Q��S\ &�k&L�b+�+^l���,5y����������8?�ΉM��
�Ū���|�blY+��{Aʑ">����{�DX��r�t��B�N}��W\J�vT�%�� �Di�����{J����[��v�֩���8c�J'�\kT�����GDͦ�ȓ&^r�!�;���R7�Z*�x�=���2i+��vb���.<���p8x�R@uۄ�Di�Y��<�`���;�I�|�xhdL����5=�7w��O��R� �Փ�&(���z2>���f��#Ml_�Ѱ�������D#�S�y�J�kq���dDZ6��.t��ox���t�K6J��Dy���c�
,6��0x���/Q�z��kMlo6I�F+�I��|�8cu�&�M}j-�����T�0��d��%0Ŭc�W�6��3��	TX)��  *S��!��NE�!dL�ˋ5�ӱǗ��}(q&�H�u-�Vb��V��ԩɫd�ںU!1�	5��3Q�Ǿ�kj�ӵ�H	�R�47���t��� ^_��:��0u�2��$xZ����%���(�_���$��v+��ei��4K:�}պ�ڜ�Wr}�1�=_#�>�_�f���Ì�B�.�m�"nsh�SF��|�L
�ĊЄ��+8�i ��������6�	�8�� έW�4iN|r�ҔuX��L,���i�������W��k�ڄ(��$in7w��xY��1�u?!�Jh�Ԯ�q��.�(O�DB7���,.N�o���I�R��@E]0�<t�3���&ܫ�T[$�HA�^A���8J�HR����Ka�DuX>O�<����V	�[�I�:b9f/с�Ո'V�r����ά�-��V[�D�,�Ѷ2z� P_m�_��L�(/��%W�����_0{$dǕ��^\L
6F��h�աcɷ�g��ߗ���~69��P
�1�_q�#���o��M�$<6��)���+d0�����Q%�1����庬(�R��8�W;�b%7Ay{�|忮����$�{��AZ�z\ b�;���бq�y�?�v�9j�͂�`�Z�1�MvY�����'�b:ۇLV�����t�^��1�y�#�a�� �z|���6]�����W��e
��a��v�bb�T��n,�HZ�WS�
u&�њ��c�q��=�C�xv+$=y��Ľ#ڞ�9�	�^X0�4l�g�S�yh��y?�`"��AH�!Aj�n�΍6^I�5�
U4#E��P��`?^ӈ�7'������,z�����5�N��O�f}�!����&����E�}r=rD��JLlӟ+�����a���v"|��1HX�bF`Cl����u�Ds=�3�{�'���	*g���7w�A�߽x��=zc]���%.��a,��]����)�x:)�-[���R���Xz��9�;vqTW�V}	�@\��i��s�
Ff+V�,��.�#��D6��뫪r�~�6��=bE.wȵ:~����D1<@��N��u�<,�QZV�n\�`��,�Sh�d�nqF��C��A�=���c�����y$J��X���_���!��eefD�E;x
�g��|��X�޽�������GlR ���9�p���)L &�S1E��P���3r3��`��9mĵ��ҹ��~������d3�]!+�-��W5/?%�l�����[��h�����[{�ʊ�0t�9~4�����9O4�M�w��
#6m-8?\X����9 O�����ÿoT�m�H�s�nr�O9��D���)�˯Ed�R�)t���G���y&��&��$�E�Ei^�n V���R����)��Z�1�㕂�y7]�J�*�#���	[w�1-�$���S�Tt!7Qϸ��WdUb�E,�$��[k�m~����6>�������T �l���?m�����rU��j��n�4�a�Lá�4��G	�}�k�M �	�(�f�ޔ�&FQ��҉监�d�a�[�#�GE^:��+�-o,���dM=�M��� �v�!i9�TUc�0¬6�_�������ȾJJzrS�J<��^�Z��kx�� w��S>&�⸰L�>DY��l%f���&k��h���+����nXF�6
��S����Wy�@u�-�\x�`U�y��C�A���Ӆ������� �}s��c��^���*�A���>���	��C:�,�I���r���To�QMrX�=UܵL�*���f���ъ���7ݒ�J�rf���z����Z�>�{!ϩ=�(?p(�L��ow�Ƞ�ت�Ƈ�*��� _��k��+�\F���L�{?��H�f�?�
w
�Pz��95@Y��˜fyF�xG��#A���4;[suť��ݤ!�NW��&�])c� {�t���8�!��yG&0��0�ЌámU�%�:��!���P,٦u	�>1u?�ߒ�5^j�p�s���j9	��ug�(�y��F,�7����|�{���\{2�R�� ��lT�v.���]���<�5�}`��YB���q��&@(o�w�cv����%")� �Ν���Z�x�Ȳ�'m<��?��]D/K�|e�$լ�t\XH�X���6�Ԇb&�v���3���y��2{I����4"Zf�����)�y���ɘ�R�A���4�S���RO�7m�����ŦmP^�c�f�ީ0��u��'T(8
:������]���_d����@Ľz���pő d�JU'y���Bᵿi�:mTgIZ�PirV!=~�������D�'�s�'D�I8�X�u�}+F_Y-��G�?4���kz�-�����fa�~�����4�6	�{��dG���l��:�( �p��\�#g�7�s�d��j'����UCc��;�Y��WFE���4P�y��,���8��r���> ��p Be�i}w%u9 ~Sf�h ͊�,��D�'_Ֆ�]���]a�i܎�$�V�/�$���R��H\�aR`�e�xݥF����+6���W+��B�5̯Y�|�!���W�6�{�C�Y��j^��	'(�����Úͩ��R��o�U�k��W�X��#J��.k}�_3"�/y$�� �f����%x������d�\����_���t#@<�jc��J+�[YBq�Wo����D���F{U���M��	A`VXi�{j�Ԑ�t����mx׸v�����]g��y����Y�5ɑs�p�� ț��D�%��wn�@�U��
���:f3�q�c�}$�Mo.YI���1�}N|I��������P"�㈼�)���!��Hv�6�Z�ZJ������x
o��&.f�`�M����ta�nx��-e%��%f�%w�bw�3O#:7yȤi�.�� �!	��k)�)`���;��
30c	�g��-�阮h=���0��4�%v'��6z��������L���<p�@����& $l:&���L�(�_̧ ���@���Z̫��`�A���U��Q
H|n;�l���N��iŵ&���-�nt�4���Ӂn�n�{'�ń�Ǧ�,g��Vh�����O��`&��I̔�jF��5�n�<�lCn�Zd}Z\b�[��T�a'aok��ɟ�n=M����������]%��rC-�	��Kl��?p:��KAyG�T��G�,{G��{Q��\m�-����%�0�W�C����[u�:����C�W=I��U�(1vu�����W�}�ۙ�J>�|W-#��`���s"�?���P�ݹ����
~S���{Qjg��6��ƋX`uO����9+2�A��2�	��p����O?����tC��_K��@���"���}�bcO�A��~����wH�|��0�(��r\�&A7:����\	8Z�!I�^Ǿ�Q}i��K쵪�Kʣ�1|8��?_V,h�Ս8���L1숅�GC;t���i�J^b����/��k����E�[\s<��o*�y�Xm�q��(�@>�,5^��"�k�k,vce��U�T����/̊�b��@�g��5�f�o�N��/a��q~�&�o*��̑����0e~x:/�����˖�;����4A�Im��C�$s���~Y��>�^k=Ѐ�@�;�Iٹ"f�z&7�+������XrP<�� �ܱy,S���0��M���19����
�T�L� �� @������M�X/���(uu��X���8M�Ű|�v��8���D+�vؓbEA 0k�%�{���\q�(VDc���쮝�ՠ�oMw��"v�Ƅ�1Ԑs-^A�
]
�� �h�XT�݃�^�'��q��.IY1��RV�	��
�Ȇ�-QK�j���e�aDT5=^W>�H����r$ͱc���ov�2_�W|P)�"	w����;��x�q�[�U�s u��y�������c����7�еv_���&�F��{���̄Q��ɇvA��!`f�M�z5��LL����I��'�t�MU�{@:�I(&�D�`��aU���ʌ���h�`�1����t�$Y�*��N�c��(?e�A.8�s�|�KAG�����b�����	�.�)T�6���W���!�TA?���u�r��fP�y~�i��R�i��? �_���멠�6���|��[-��� $U�\ѹ$�f��������n�K������˼����>$?�y*u঵�O�r��E�G�*yȁ3ɖ-tc-�0�I�W�B�1<�1^mV�����Ҏ��FB$ڇ����M�c�a-FLE��%FB|�C����vB�؛Ƙ�κW�x�*U�v��zJu��S�?u$=u�D�h�t��k#%��08�G9��r�ĺ3�o�B�A�^l�C�� *]�����F��V�y�I�EU��,�i
T�7��#�rL��ڑ;�Ҭ���r��"�T�E<�����H��	b"��υ�`�$)�۔ù4�X|����5��0O�������F���ԘEUו:$����Z����H�����9�1a�T��_��?+l�����/�:��[�cD-Tr�2V�|���,Q��l�o���\Q>Tb�kt���ҳ�i��Z��A��'ȣB`�KH����y���'
�xg�
E�����Yҩ���ؙ�跞ŗ"����y� ��Z��ӑ �2]�,U*[g(�����[���y3 �D�Q�Jix-�ݹ�6������;TD���\�
jb��i-�3L��.s��_CMb+����~���qQ��[L�Nw�'S$�d���QfWMT�J-Ƚ=��A ���L� �g��!�t�C�ZC�2U�M	u8�y�t�;͇�iIh�:�]A�F7�Ђ�F���!�(����#��e���S�2C�������hB���F��>uRd����/�6w9
E���/��ھ��35 �����1iQɌ���2~�k����3/y;j�U����ӖXuPV�R�)��ʖ�<"Z#U���9q`?:ahzO�;aJ2Y�pC�c���U��o�j�u��EU����*`!��J�ʸы��!���@�_)�ՙ��`��T�y!OMa�o���}Y�DI�	�E���7z]n�EV��K�(~�8��%�}
���F�3]�ۛ��;�16=%�M�B>]:x���'K:�HE��4M�Ճ����2�N!�h3��^���6샀��D���/�E+�"��.c0C��|�2�a\��چ �Ōs������5sH-Dt���!Ķ� 8�e�a,ˡ[S�4N�B�=��u���a�aM�K;�7M�i.�XW��r���|�t<�U�`M,�Z�����y��#��u�2��J�0�GÙ���n�ݺ�5���"��IQ�k�tVس�a�I;%1�8�Wl[����_-����c��=3���'�:�b�S,wɿ��g�����GH�Y�_���T4�ų�"F[�ޑ�K�5�B�ȿ�i���%`��l-h�B!i?f�/xu_/G�&��+^�bJ��F�2�~Zj��6���)�u.6�w^�ϼ,�9�Q2��<�]9C�D9Dd8$e�Cf��z�rd'rC\�'c��I�)GPi� ��_��A�}�78�5��'�³��n�Ӏ^X=D(�?��W�l��E��u0�,�VK�^��Rxt]���l�F�@g`CmҺ��Wݞ�	TB	�'R��ڻ�0r��U�G+0H�����b.��r$y�]{�gu� �R��L�OX�0kswfB-�)L�����<f912�0�De���:�N$�d����zDf�([���e,c���Ē{-$�Ǻ�%o�8{�ď('��N�{p�z��>I���I%$��D"�w ���gN���f�2�2&��ۛY�ձ<�]�����.taDs�Ωr�C�(�#�&�o7N!	����W�_�KvTM��~���yq����U�K�b� ��KN��4�H*[��grx夝����	-s/li�lkC�E��^��"'pJ'��HJ�6�Y�D9���4��p�v��,|ʙ�9����+ay����E���0~���3�d�i@z|�ɛ�������$y|���l`0�9A��
���d�N��%_����?�����(�c�C8|J.j��O� �2�GG�;��=�*^,Ev�~��O[�S4B�.7������
[NTPǐ��i�Ѷ�~�[+?��~���k\�u�<|�0����Ң���#����?�iI�|jR�aϹ?��� �=����e�j)�T�v�EE)��:�����ݛY��v�n"��<FILz!Ca��H����>��*n��u��c��,_���C.���j���m����Q�̮�ІV���~O�:;��~��Q�b��G�|�Z�/"�=���3D�?���&�Mq͒ˡ���2(��xJ#eWĒ�V�OأɌ�#탈?|��um�Ł��3�����Uz�q��F�U�|�]�&��;�LtK����_*��5<J{�;�3��z7�bv�,u^Q#�Ń6��!:�������}}��b����C���9`<;�EyN�6
u�6�uy�w�ϻ�c��2#��'��&,��z|�OR��=)��i+b��iΈC$��5ņ��F�ìiNjs�(����L[,��6+W{�:�b��h��'�ށ�I�bo{����J
���A���0D��:�y�ǓT�z���� y0�w���dYs������d��u�g�KI�6!;���o���Ӡ��m��\O�	��>@�����+G�{��Ii	�4Ij�D��@^��us%N�#�u��G�ǂ-��v���U)�����rA#×�gFq�KC���7���`'�j�-g2(#��3<���<�zO��ƥ�8b��}0kI,̰/�o�s��3^v!*�P`P�=��\*].��Z�/T���,Z��~»/x�k�� �#hԆ�Q�t�&V�x~���u�e��ه����{��ԡ�?'�9�Hù)P�������e����$[���Iq-u���7��2�d�+�]��YE��'�N�hmjC~���ˣz�'U�[�yr?9�Cʪ��"�@�k8vÐu��W0Kmgk�j������I���m��92�ҵTbǏI��tٻ ��ܸ��|�E\����R�ԛ5�;�gz�;��[{-��;zT�X�A`�V����8�h�f�^@?�/s&v���b�nqR���
 o#T^��Y��!�4��#��b)N4B��}�fg�!ؠ���6S�cT6\"����Կ���F���Č?
���>3=�y��௢�',�~���$��M!�|�;$���/�y��9�Tv�4����	|U��Tr�C��|�P^��\�*��yet���[կ�0�9|�%��X���w�r�k�نyԲkR�D��ZtF߲IEz�Eq�px!���"��J��!�}9/Rjs��{'3�)K����0���2g">F�=p&b���Ec?��Խ �B=����V�ۗntK5�ߖԩ��tYly����_��=��c��D�b�/���aC��Q��T[L�K-�u�$�3�D�;mJ�:�;tĆˮ^�,_���&�M#�rq��80xVV�	w7�]�����F�Ό�N�������w%{�XfC��H��J�r�&$��q;�4`W6I�h���kX��Қ���;��ke�7�#�M?G�N �
�9�縵.aE��yO��7���8���Y�
*%��;CF~�1�,���)�����|uu5)�>_�؍�&f{`Kr43G�J�~���{d�<7����uô
A���������9#���w8��W�8*�_�HͪVZ��	����.��+3$�d%� �O���D>�6r�)��:��Q1a�&��֟���X��&��7���}+<�c�m�mP�Ӻ`Vq}��R0C}(�SLB!���,O��I4��?�TV������N_����������#�)|�/X���g梕S�mzU�zZCƸ���Ƅ��E���b�	�s�"�+�@����~/�����d�ii ���gC�wM^��1q(�s��YWy���Ɋ�Io��F5�ޑ.�|��(��i�c��d�����&�(\�e�
��k�7FOUzӂQ��_�O�;��8�`��7���g����T��i��i9sݖcD����LlfՁ|�����G?��O�S�~/xA;��O���'�z$P�y_PN2s���I�]�<�/Z#tr��v_�!I!�lp���x�����i�EWn���%UR_�����z�8�;9��5��5�1�h䊖O��S��頳8����L����KRt�~��J�{� ����H���ϲ�(���8VD	�o1"mפnw�}��ߊ��k�z�M���#<��ZN<Ty�(In���tK<��I&����J��ɨr�S �M��Nf#H�Ԋ9,p��x	�cB��L?��o�^�����0��n�6/���J�& sa@�	��1 ����v]��D����93F#z{���k�2��i��I��M�z9���&o�����V����?$����=�>�*�!7a�ROG{1�k�}z�6�o����X]�;Ӝ꾙��ȁE��6���zz��Q�BR046�3�|�;�C�m�o��]�����+�������rm�N>�Z�ʯ&�����!a./LUr�Y#�5��ic*��Θ���g�g*5�M5�z���H���~��������u�8Lm�ܰ2:q�ElXMO��FGm}�af߱Y59���b���j=��cr�0M�J9@��8�x��U��}���[gv[D�������҂t��	V�Z��T��6A�O���zڪ훚�~��d�*����A%,����W3��:��r$�	��YV�)��~|K�>��U	$�3��٬�LEn�<��O�����8E�DOi��Bh���A����_�
��j��h���������+��t�-N�J揉;$�b�ښ�8{�B�I��Ǽ�HI�0�'�=�"��\��)�iK6����P��l[o���:c�cy��N?A�G���Ғa�C��y\�=��g��0�l�������0�($�gY9�GʋR�½4M��7��r�B2�цM�p�\������	��z�GM��[)N��Q~����u�x0�lh���2�ʬy� V�2�?7�&/~��1@ ��]���+ 5�2X>0>��z9{������������N˸0����U�Sg����P7��_y�t���7��XP~ ��o�gjoQ_����{́ӫ�����F!�ö�Rǖ����՝��TJ���;�#���kW;S��X�M`� �ŏ7��!��HV���6�{.$v?y/cYM���L5�p>Y�*DX�1�P�K����VzE��YU���A�,t��p�(H�<�TfQI��Ă(�h���`J_S]�L�-,@�X-0y���mmS�S��sտm������iʐnF����B���D��.��i#ɼ�����>s�L�[	@S<�ثA�؟��%	 4M�~Y��t��Z����|�@�sp�Qz��*�kdf����k��&0"�6�1�(�_���� �@<Nc�3皋��p��%3�z/��$�f�w�?yV�*�3�A�+�)z��r��Nܞ�nd;�JcQŀB�w�ҍG �r����m�l��5�<G�1#q(j�T�(���6�TL¼��q!~�EZ3vt��:��-� �\�e�a�H(ئ���@Ջ���m8 ]��Ί��u:u���㉱�b⯍ ʼ�J�\;,N���b��c�������b�rڲ5%�]�\�bD�����������x"����I���r��yFz��-�Q�K�r=q+�ǒ �>�*������թ6�p|?X�:�.=U��׈��q�7:{s��7�Ҍ�ZB.e+��hJʵ��ݸ��u��mbZ�l}��ɷ0�?w��{���&��ZFq��M.¯���z�Z��=y(��Z	Y��Fo$�=�\��=Vp�d��
�6Gd��!���(~lqN^?��+؄*L�e��(~��u��9-��o!���[���Yna	�(���:��Q�O�����-���;��g.áǨ�Zǃ��>���Q�T�L?[e�sc���2�v���ok'g���]d:�sz�O�)҃,;)�t�U�Q�"ә���+�}�y��E})�DZ���V�Hl�MSA����-���=r7R���R#\��cgģX^�6A';���L"�k� �D �&��|�s�d�qa@t��2[7x)��dChg2?�	��6>#kb������Ȧ�jʛ(K�m%�:Ɏ.'T���c!"�N[;����:p\{@�Ͷ��gs��e6Q�?*)H��?R�{ZncsP\��~3Gz8 ��j����X"g�c9wM�H�;Q��>��]��݂~��PE.�X5��6�`������+Ґp�����y�wk�.�5G�9x�+����J2�@<�߭L�X���	XӢ�""c@����h]GS�m`a���,�3�8�EIs�R"wa1��|Nu�I*��[���.�?��)��Oe+�_Ə>p$�M�>e�Ȋg+�*vպ�H�;s�S�5Jd�U�OpD�ƫ
i؝�k璤{ɇ���(�����QT�`L�:�a��daǻrDp��}�)]35�GA: D�R���c��R�	�)Ж�S�&<e�\����H����}���^��
n�EN��g ��v�A4�n�	��d�2,���2{zU������<K���2�p��[C�h:��La���!F�V8L���L��r�P4������V��R�޵LeĔ�p�UL���S�ۇ�V��/���)>	���xqMqL��)J�`��H�G����)$W�ܝZ�>���!�@��P����y��}��b���`	���:4�Wiv(7.2_c�[A$�ݥ�*K���
��)�a�^N>A�$�����|�b8s ?fM�zR���޴�$5��"n��ۘf�1�h���J�2T��BTq���_ҡ�t��n�v������O�����ʉ���dT�Xz�;�}su��W��=��u5f�����V�� h�u������|-н&�'각����&W��/��i��/NږKJ�;&�#Ds(��S�h5%�62���a)�9!ëL�����,+e"ANg���*LCU\��.`H��8���J��n��&�O0�/��X���v�l�":�sZ��Ä	}�QӪ���HA,&�w�</��U��JM(e����/}��c�n�D�k���G�m��oWk����a5:�s�B�5����_׺4���)b�����k�����}c�@�y�PSFD)�uQVp&���{KA�b�����$o �g��{+�5ڱR��X���Ad�%e�J�d�9L��&bM9�)�e��O'׌2*d�A�Q.�v�;O��?��n����Qj\)���O�;M�͈r�hWu.���9-+��q���&��쿣8X�·ou�ek�S͂l�i�=�ȏ���BXJ�ѓ6�ԵU��ԫx1��`�<�������񦪼��^���uᦠ��j��W��T-�`�@6 	�1�L�qAy	'<'@!��v�
]��)��Oe���� ���c�Y@��Q5�O
�-Q�yn��[f�]i'����Lt�OS�F���{� Q+ۣ�b��c\O�����r0p6�>?N1�O���}H2��+;<2��.;fQ��.�15sH.�B�&�*I/�1�A��Ɯr-�K��|qm�O�����ul���U@�)�yԵI�?Ezg��,ɖ��
a�wl�����=O/���'m,�T� ��O���p<Ayɣ?�f��R���<60��GtAӡ�	k�
�{��,�����cF�h�����ȫ����-�k[���$� ��F=�<׌�����]�畗Ϟ7*��P�^�^�.�4��i�|r��R����k����_3�h�	$�北\7�`ä���j-��8�y P�r2�˰�v6�V#�Լ�� �-S�>H#�;���:w���O�ɾ�|	b�G/�n�r�lR6���L��.1����5�&S�آ�S�%Җ|p=uT��$��~Զ���;�b��?fE<a��5�t��8~=|\^��.vP�I��'����3�xBk��r	"���?b%[ɡt!�26�[�x�O�\=�{��ée�W��<�ʚ�~m[r|�g�b�@a�<���n{���(V��$��똵U�?��'�С�z`�M' �����p���X���zJDHGwu (�d	Yy�+���<��
�����0D��1ւ��u?�T��/�J�xd�1	y���M�D��k��;&LR �9�Իf�2/O|�Q�T���W͗=�����Ɲ�他��B�O.���X��˸o�f ;#�A��f#�qϛ�>
x[=����}lDv�/�BwG��u����عG	 |�������NOp�Ztq�J�5���[�.!��C��}�����A�.�Jϴny�}�sX1J���X�$����z��[� �K,#���Yg���A�n���u����F{�횸�*���0�a������i���XI���:@�N��:��3�TU�P:�͎i��'.�1t���#B�(�2�}C��`�/�
KtVe��� fE� ���M@+gm���X��Sg׺���Ј���-�tƒT���7�@�%iE]z��0z»�"b;ڛl�4�'*���n�i���-a�E�I}V�ʋ��J�_�)S�;aT����?�y�=�a%%����w��j\�����$�A��W\��D$�
li6�jv���t|m�$:»�lI*X�f�I6�ո���M��,_pF�H�@�,�����M]uq$s���7���"�[o1�f~#tb�Z�u��U��'Y�݀���Y�0�a��j�-�
S�S��s�o�4`�]2������d.��V;�,���I �KTKE&r�i�]$�mc�hS��7�t�H
;�A���,��c�� ����� �~9N8dJ>m��#-Z������;���P,�>�s-������Ji��/�l�[��0�����X��/WP��@���?Z&�Oh���Ţ	΅�Vh��2��3w/`�V�nG��
f��c�B�ف	�?�#g8�l��_�^�xxQ���$#5��D�
��Y�L	8[������'N���M��ǖ+�!� �;E�
�76���}HqT3�5[&闧chi? ̀�e޴d�,�5�s���˳3:}rQ
#X���b��ȋ�a +���|�Z?�n��fm�_gD��?w4�D�=(�Q��P�d;�r�0R �ax\Έ��� h�Ñ�%���Q1�wܗ�E�MD?����q'cjh{���	�j�X�t-��<�Gr�o�I:O�J�KKZ,C�DgdYx�LE@5�	������Y:!T��^���U�����G��]����-���g��
��b@�	�:���$������ق�j-�d�y<y��/�I㨄X�7�-�������»�=���J��Q\� �:z)����kG�}��?+���;C6:9����;;�ѭ@(���b���z��,�L��a����\q�4$Ϣd�;�׿��/�,�Q��vJJ��<�9:-5�ĨI�=�Q�$C��I�(i�x\Ѹլ��j�(I1��/�;�/^�$��_�O��B�Q����=neîP��IY��\0 �� �6B��1\�|��;?�q����~����˓�E���&Z�$�gY=���� �},�!��|���M��YLL�.2�=����X�(��
gS�^#�(����٣m�6ov�7���̈́��
�g�P��\&�������t�:�Dշ�r�J%Lta;0�9��&7�0���ߍ��	�����5/���~�肋�����ˏ��^4!�鳒�%7!.p�a�.&���3�M��G[Y�cM�T� ���:������z�=�s�b��qF�b�c�/��$\��> �هT�5���:	����/�d>��G6{ql��B��\]�msL��2d�d�&�����9�y�֬�k=�{P去O�If�Ή|f�6^�!����fZ�S,����sm��5r%�>ܵ�xˏ4��G�%�(� �T2����7�c�"�_�9JF�L���}i9Uq-.��"d��L}�ِ��ǂ,���'#W�ʉ@h�4�2=vt��J�Cj7-��!�v	P�,��V��3�u�U�&'�\o�ۻG~v�s5�* nߟQ| W��h��4 ��.�OUK���8cTL���@�I���oxb��J.�J	KU�w$n�ƑV��fD͓M�^�Y��Q`��vk��dn@BF8���B����H��y�T�i]��?4Zui��	2=�~��� �-l�H���Dx�]����������l$H��sB�Ͽ7׮e"��_�o_�#l͞syY�N��i/�*"m�����
���+�mI�x�-�����\��̇�� �1�j'ʪ�ŉ�� �asuF�]�Ot�5i»^}yu�]�
M�٫li�f%n���8�o���
�,\7(�2d]���&7�	�����0PGǕd������^%��MB��H[�Ȉ��������C2i8��M�6BX.".)>��1d'֌��3c�Ҹ	��l�L�(4��v߶|2��L�Z�O��� GV��c+�Gf(K"?�����LƐM�]�葧t�Nd�b�f��F�]oB?�&�芝�Ko�+?c����0X��
�C׸�7�x�vWQJk_K��u?؋�Tٔo����P��m>7W���)d����u�7��|�ݺ�J$^��^�D�}�ߒb�ÃDŎ�6�Ƒ̐ ,��~��ev^����_K�����<K�`��ߓ�Hv��g��A�ԑ��ڇ?.M�e)\��'Ui1��Q[!%����I�D�\w��#)Q���k��_�ra��bg�!#]���Z�M�����!���]YB��W�- �gxՆ�.�,~!����D���b_��L"��%X~�lg�.�-ho��)�Cp�m�b��h�"R�QC7���-W���@иڟ&�nB��)��iM��/& 2�u�Z ���-�΍���/"�<r�N�ˆ4��K<�Pm�7�&鷥q�6�2,}F��36�s�D�l�?�n�����뒝t�&���T�Nҟ�S�d��/��Ql^�N��{f���t���Q
�2�:,�+���4�tp�֍�����6�m�2�\��$�Ray��G��U�H`�j�C�!�Փ�����/&�B�c��&^R1/<�#�bʉp�^�;�����t�`��C�}�.N�̒29���b���K���b�Ï�2��fY�P��eI�v;��L�p�z��Fp��æ6�%����7���T	���;iRxc3<�S݋ci�h��pv�y��������'��Q���@�dN,�O�6=���Cen,D΂�.�!����)HIx0y�F 4���5Oe$�g�Q����#q�fPM�ZR~"Cy.`�褰�k)�W�V�³���eˠ>N�6{�[�9�a+]`b�������'��;zATK�I�\��w6E[��C����}������|����?.s��y���3�|�6ǭv�lq�B?�bX�z��ˆ�p��AO�,�_ �acLa���,�� ym��erˏ������Q5Շ�b,�)�VT��e�Xvu-{�� �H�	�v���hg�|��n��5�`�Mo�w]i8xY*�՚��6��v�bxR[�q�:H��tsto��M�PF�#?�RRW�����!N"��O����w�j�Q#��UZe �1���7Gn��CN�� �KL����T�+�Y��5�2 .e����$�°s0�����0X�h	��>�I��&�<DV�B�F�C�/t���}E�0U�s�Y9xX a��S�� cx݂@I~_��΢/����Ʊ�;���;�k���63U�V~S�/�T��$��7����H�h11�%e�'�2V�|���@������~�r��T�՝���Q��;,�F5����w1>U�H��,l�_�<�;�,�A��k�ٸ�j���r�b(p-H�ڕ+=!�4��?@�G3����z�M|'o���oO�N-��;G�`�����9&�r/$K�gL�=�]0�j!�sI.[$$��uKK���3��b������|�������p[<�O�W� �0�9�:Q�k�Kr�9G��B$�pcR���jC�0��2Di�jx�f0?ա�N�#�L��=�J��a����z݈5�&o�a����	K��I�#����6���0��B�-��4�t�ͬ	Q=m��$/�:��Tz�^V�U'�[T%������0��a�n�*מc���?C:���as�X#�;.�.x�}�������@L��s��M���u�$���#��e6D>�4��o�DF���2�5�����ͬKT���͎�VM���sq��od�6|��+:ͺ�����}!D�b;����#��w����m�p n+�\�4ma���ٰ�;�s�ʙ��}
+`��5�8�X@�9ag�st���C��0�]���_��YD�W��@�6���vXͰ�3Vqnґ�(�h�R�=C,,��k�k|T��GU�Q~�uasE=�&����	>B'e�vM�b����S� 	0�\����ۧ�����M(D�y�d(+�1���7B+*������5ר�����t���}�C�<�,��_�����wAv͖s
N�q�7`��~�0h;ې�h��D���P.��浊j���g)�G4���`�}X�em�w��Cl���d��\Evr��Z�U�Ǟ�0�'{�s�^��-���a����;��zi8�;u��D����
��KZY#֪G��SD�;-pH��0�>�^Dq"�c�Y=��;xnZ'�⼀�[}M�����ɥ#%�oG:^�M�j��9�(�Q�&+y���\9���<����$7QЌ��5Z�Njc1��_S����Q�~&ul�����}���%��_�8�A�$u%m+�?썣��#Z�gM��#T��e���K41ag�*6Ȟ"�^��Y�1Iu���G���s��Bk�)r��8�ZT m2Gw�t����|.0�ʦ4d6;l��%�g��ma{E�w+�5������n���zM��P�~s�<�������aJ߸��q_ރ�<�k�f%�o<44�?�Y̫ĥjH9�z2$��'���b����2>8���:��:.E������X�������8�L������:���vv�7 q��� y���P��I�Z���!�S��\{���[�`?�z�h���-��JQ��#L���!b��:�1�DD�Τ-!P/,�^�)�{�1q�Gt\����Y�T۟�i�KqG�G�/n���N�YV��_̡Zx���;M����Z���n2- ���mo�$�����/�`;��+d�I�(�&�(����]W���\1M������
�Y,���M��إs�G(�g���� 6 ��m��7�D��Gf���о��"�R&@�GK����x�����%m#�?=)�K�l�5?�4]�&�y�_3�&�V��T;���L-�%����q�4<�=ʢ^����7U]zm6����wRe��3
0_��q?X�\C����AX�Y�Y��8���F)�iz�|/��������P:�� �]D�#u@2��}.�C��X����$�k\J�v�pFA#�zDE�Ȇ?W6k7=m} ��Kչ9�-�@ւ~�~�p�x��vA�#0o�-`�B�b��PCˇ�(���lc������A�М���S7�0<b=s�G��sT d��Yl�C�R��i�.�˫�ѧl�T#�;�t��u銎i�/s�F<c�eTj#�� ڬ��PG߱/�*#+���E���v���I���~~%��F��aZ�{�紤4��B�(�[��8?� 6���*er�����2�`w����V�N��Ʋv�BEY�BJ���Fg�.�����y�*J2Al{��y5�Bc������ϳ�f�N�ZK��f�p����T�}�^��#y��I_��Dl�;V�[X�>/n�<����h��q��hUl5.,��'��S�!fw,��Y�3�-�5_�a���Ðnu��OG�}6����j$mάl܀$.O��Xn+�>0^O��#ui�Yu!:z���L��n�A������\�2�L֕"�Q�=��"a4~[���J�����$
3�$k*�i�0cRn��,�Dfc�r��I'�w�HB�A�6익�����U W�äC
xE�5���Զ͑+��)�h
X���+�z��}5��՛��<H2{]hY�EkG5����u�:�3P&'S�ԕ��3�}0Oe�t���ࣰQE�����w��_�4�#�u���=F�a5�]����7��X���մ�X-Ԧ��w*o�g�#e����mg��KQ�~����%g
��<��{�k��-�?���4����[C��>+B��҄r�S�{���o�X4�`��6��ʖ��ˊc������@���8�w���B	D8f�t��_r�9����R<ρ��<�~Y)��=�~O�lS|ek���V�R�_��gmw�P���o-{���EHSJS8��2�x85�f �F�L]���	�$���
�ɯ�>�w�0U�!f�=,*Qn洃�j�G�޲g�|�\Z��X�|�X�sׯ��Xw	U�ҡ)
�ǂw�a𾍏Ȱt�)}��䵬�^<r.[�t��9%�j��rs<���/�Y\�_ �RJb6#(-�j$������`�u�繳r�$���C'�|�>�2��#�H�K���/��1Ӵ��?w�Ft��)"n�eyU��W�Z*�w�%P��:���.�˒{�'`�F�ÒxC�$��� �T��}��"!3퐲�*��|��-��L�sX���ل]h�]���?�l�g�2	��h�ˁF0�]4��@�x�2M{� +_�b����ێ�fK"�>X�~dS�0f�?-f���Ij�(E�{g��]mި���[���By?&4Á}�>+%��e�Ol2����Q�^���?�Ptg�T�B�N����/::M�g�a����i�O���������s�&��x�{���6������T������s�Od��b�L�f�_�7VO߲oN�/%_𥳐��Rl��^�����I���ݮ7#I�UC��4�X�XA�U5fbb��ڲ�]������bq �kkW:CKg�W��%3q�����?%+X��'�����=g-D�l(C|#�Sb�8lUj@� �]s���[�k�ʺt?HFJ�Q�v�P-�;�쁍����b0�j���ކ�@O�wFE:e�b���m̀�}��,�8����Y�tK�"ˠ�B���赡��>Ս�u�� ��9��u䕯��c�2��v0�H{xeA�g_8�*�JE��)F��1C���!"%D�hϦ�jf�6��I[��̈�y2Wr�?���6���z�j�����GD �,=} �i�*Vޱ�B�Z. ��P6�����F�驕�N��`[��{vGk>�*!�w`NO�Nf�u�%9��]�>�wj�b�ʒ�y ��ǐSz�M�/׃)]�6���C�-�&�G󩒎��d�Y�A D�ޤ�{����M��6�MV�q:O�H��.��w�ΨIs{@m�� �K��4���{=x���r�����*B'R�$��Y/��|��Kh�.�QnRBs�rb���f�I��P���o)ң/Oq��˄�<��θ	W/`"t�����\��Z\p,[��>��@p���-�ѯD�'>@w34���h��_�Qe��2U��IکTZ���s��l���C�u�W����!��U(�x܋k�(�&(�Lآ��~�����l�K=�~e���\��G$��Gp���ZT��fgVgӜZ(WIe�ѩ��W���p̓�z-G_��)an�0�ɖ�x��u��u�1�Ȏ+��W��{�z\�ED��J���X�0�}���]XSv��
Ѧ:�jq���r\d�K�hU�2�(7y�:ћ��o'�`.M�>�S��#yl��_TL��xɻ9���6��E��rz���U��t�U�,��l�`�N����K��1�Vh��}�� �	c���2}�G����1���;�]	�(+Q	;�*dT�U�m+���xX���$���=���Z_�%oe����q�|(�+є�@H�xsww��F�_��r�N�T5b�#��Wh�?x��K��St��󡤰�L�,%Ompi�P��l�y�3�6���գJ&<�($�s�:�`��Am��p3�	�z��s���'V���
�^R������:�µ����n����9�'�%[Ds�p��t/�/D��)����r;kD
�4�����uڕi/>@��A����9���J)0�AZ~�m�����
�<�A���^U/��5���E�3�P$	YiѸ�Q��Z��w�nKZ�!:4�م��z��J��EF�Jj>�#D��좃!��J�b5 �nzH���N'�X^}/�
��4�0gޱ%^���������韈e jkWL�G���@/�{�@H�2�u��*���-�O��h�m��1]�7��<>�_���G�Լ�q��r�!t2 m���E���}+�Ũ��I�	�t��t2a?'���)e�y$�T/��k����s}lV8�v�AR�ae����C�ѥK�]璯t#�=yt-�#Lˠ�W%�C�mI�D���C{�_}�b���ˤ7�$��q���ni��B�-F{ ���,8B��f/%?Op�/�P��ȘCu�W��\��������\D�8��}�$�,�:L��f�j��â���j��x|cnǘED�^�����P�xG�y�L|���a��Q�9i��=�*Nm���T���ڮA��.3x�LB8��������&�7�$�tq	�G{�!���B��84}��?�n���*���։?�c�n�c�߆M`b�&�5�`��4K6�L���Q_�	,�Z�/�I�2*i=٥�x �w!�ޠ�4Z^9t�p砅kw' �t�M?�SmbC�	�$�U����w�tbUvYBfx1����6���낽"Y���ਣX�i�fq�_�cTSF�գ-]a�)�q���Zei���Zޭ��O�S	��]U�'Y�i�e_П�y~`�W��35�nX���ߴůT4j��kqo�X�}���L��S��l�fd6<$1�nᮩ�z�#���������5s�Qf�BJ��a3�:���'	ϯV���y�L����<�M�K�K���d�'4����{�k���T������v��#��2p.|0�|7#�W��ː:�6�|��u��ܙ���1�g��O��F����r�h1��^�Ϟ�� <l�4���O�y�5]�a�>sa+F�:����,ǐuf���y�G}��"�%\)�'���;x6�=�?w)������m)Ī��К&Z;���nr��t(��|Eһ�(`D&dR���Z�=<�6V_=�oM�#����,�iPJC�'xF�e �N��Z3P8O����?�6\�c�[�0�R�ר$�������\he�Jnt,�":г��Te)�W!�6w��Yw
���P�ʔ�K�bǮ��5g�.+l��9K���	n��Tp O[���~evw�H�X�Wɒ��i~u>�N�Sx���l�Ϡ��]�в��79����%�+��C�TN�+��&ct*7	Ma���C�`����?pm�r[f�j(8��^O�*�u:�<:z��b~{)G�U+�S�i
#[�q,��5vvZ�V�.�/A�����`f����V��wR��H�x���/�Y
���`�:�]�wWD;����L��wl
��x�
�G�9�8a�H��|_/ü�,t����n�j��,iթQ�//���|�ІMf�rH�ӳ�q~g-��J���]� �t���ѷ��*U��8W����㯹��w$E7�]�>���}b7�4%= &���@u�1���	[����>��@W|Y�M�b��`p��җi�a����%�$��+��v%���{.j�ʆ��Y��&�t�ʧ&�~�[co��cbֽ[�����]u�S_��ޒ�hQ{Ms��;^$Zh�r�&E��=����D>D�ʉ�ۣh����S�qyE��󪊈�\S�T���2o���w�,����'S[�ąr[����4ްk�8&�p�Rg��N��u��P$�^j0�����h�Ν@�P��O��F�E�wc�6Ț�	�
���^綤:�� >�btE���gŅ�o��.͞|;:p����R��#���e��K��Nq)m���E�%��C~u��Z�e0��N��]�_��8їS!�^���emy�']��yy��w��Jh��8Wu�5a��Ȧ-0�'8��C�X�f�&#$�dz{zY�hs�]�%��0Â
�J@�}��zy?@�G���5y4д8M�m��,|ut;�\n�Ġ�~�(W�(t$ 侱 T�KŊW�o�6_��v�!ƫXoڃ��氿1�(m
Z�exT
4��"��`�u�3p@2u8��s�%m'�\|??����|���Jr]�cC]�}x��#G�̌��p���1k*;�:�{���ct5�*x<�Z!�?z+�JH��*V���I	c�[������=R1��������̾�s�3Q�9��~�hB]�{
K�Q�j�_��td��梗(1��L'�Ej��\�~�q(�gA��Q)��-��XX�9 �S%�z�Bz���d�N�9�|q��+FF��O��/Ɠ/�:�hC�[�įVgi1�����ym��u
!��R7���߶#��J�4Yl����n�/�#9N���5Cʖ����2�E}�>�	�Ŀ��!utQzJ3k��'�9��d߉��Fp�_���^�s%R�DbWF��p8Ȗo.PFh8�A�
����j����� ����?�C��Z�s�^���b���ɍ�}�iUI̸0�Y[����d��V���N���)a�a|���/�J�w�޷��������{�����P5�� �t��j��y̋b��`U�
�����FΧ�X���{�j���Θ��TT=�z�Qf��ں\�`�w�%3��O���փ�_�Q�c �ңĐ�M��4|~�d� �+�X�a�4�S��:�ǲ�߉V:CG>堲}8������uO5̘!��ۆ�#$A殎�x��Rk���h���ɧ� :s�K���Aoz�L�N/��@�X4�ܮ���"�}j���]�y���W	����v�_��(�pۈ�?��u@��y�j&^��8�C�^.�-Ű�3�	�z�x��/,�?T'���?�+�&~ʧަ᭻�q8 ]f�����k�n���}�D�
9$
F�dB��Y�Lr��TM;����n?BNAR��RkJ���7�Y�8�Z���0�b[����/^J��
cg(%���yH]��DyA����J��]`Gn�q�m�&9Ơ�aY����B��`�\v�Rd&aB��c��F4�#s��)���?!r��M����/�-Ǧ�
$y;�j+>#l9\�f��@�k�~K/�S'z�o8��u��k����<�|�b)Ko�tb�UR����Y�l�Ӄט���]���G��`޾_<�Xa�g|�{��PKu�+�w������O���U�@����%�G{���G�*v��I�e&�A��uچܵ5K-?�"�/� ���kԊ(��n&�̦��	O�*2�`�`��w�Ӳ*t̽[� ������>s&�y��n�� ��y����n�|C~�#1�<��	������a_��ZbnA�Є<F�X�i����WVd��:8sȂ��nC��M| ��#�u����c'�K�����H��p뜴9E�F��jD*(]� �*\�9)$��X�X?hD���cLь?�^g�2�%tƙ���y�G�r�j�϶�
F�5d[J7����C����Q����������������l��!=dS��#I��t�.2�����&_x�Y	�|����s�����-�D���q�cb�t|4�#���o~�h�g�V������׎wP%-ˊ�Jv�:�Ka�5�����8Y��1���Z�[���]H���L�ſ(��5�Kb���.؝��fH��-��L	����UM��<�!~V�=�Ii��)5SU���j�����[]��=��>�)����j����U��@��
q�����Ѹk2l0\���/�(��!�^����Bm�Pt�����5�sARQXe�s<(LY�XEՌĿn��C��g��>2�x�0��/�/�3'��c��A�V=��i¥�u�l\����M��,g��()~�u��i8���Ep��	��$����y8힔*&�/S��oH8�������#�<-$�lw���Ŭ"q;�x���r���":A���
E�2YN����R1Ҟ=��0J���W��yD�Ϋ(���0&B�|9&��c5j~4��	�����껜�����{+�3,Ϯ��6"�_�̭T��o�EZŜ���62Fo* iD����1���W͂U�vݎ���d���s�*Δ��8qu=�uV:��|�q&��Q;�5�ʲ8���=D�ǧ�{�"�n�`|�F
��klJ��<QLy�n��DX�c0��x\�ιք�F�YƦ���j�Z�	�H��W�:0��)�1pC�ۜ��8!�ޗ-���S�W�慃�����@�E7N�a4�i���[%�"W� ���̹&e(e|w��6��Fڰ�Q,�����$x�}0q뵏��^��4��$����/֊�[���Q��] �qh�7񞽁�k���q-������V�I�����"4���S5���K�_��i�#����O�wj�ޠ9s�կ��_P����k�����	W�6��|���C�!��8瀗JcqK�W��ѭl���$4�S(9�o*��!#y	P�� ��ck'���V����L#ГiD��:�ȓx[
G�����Y���^��,MWr8�\�({��,)W��&cx����m�JL�����;أ�<p}?�44v*F]M�
��,w�v�ɋi��ʶ�w�nۥ*����[�2����s<��i���5��S�!��t�.�K���V<�Wh9��D�{��z���F�Eߢ���3(�9oK�Cy��ۼ����R
~�L<���<]��\4v��J��I��+��yZ&*�)g��0:δ�ss9oS4�w����8P���4e[N����b�k�;Z����<C�τB���]���<�mJq@2�P��2�"Hm�2��`p��o����4�JK���4_�k�;��\����WP����B��3s�@ڢhUmT�Nb��&�Ly��ש� SGxr�2PK�0���sa�?������b�F�u�����8��nrS���j̢�ˏ�c:����z�.AC�8�Aމ@��Y��.T3�N�uUތkӒk@W���P�u���3���S�8҇JD�n|[�c|�+�-��Q4�=\�f)���k�tD%_o�l5WΦF� /@3���[X0Hq[ԓ9�V����aGc��P�]�@����E��s����k�&�s�q�=d=���.��rxw�Lϔ�]RݓY~(����ǎ���H��yn 8����PE8���7|�ۅ�<�q��UOTXԅ_(3���+#�+d�1�uW�<=1��إu�֑M+s���?�)���b�#��@���G�M�1�q�{�,������H�sT:��b�$XI�gF�#9�C����ן��4�a�� :�^����불E;�FՆ��#ډf�n�����l(Rj�J��ٌ�zZ���ʰ7��ަx\F��w뢬�
<���9�Qa��(� �,w��z��_!͹~Ӟ����N$"�L�6�s�P�q���*�W��.n~����ob�+���g�,d>��K_���A��{G������!��1��@��
bX�0�)I��dF���)��:w$�!��9���K��R/���������K���L���,���WS)������:f�-Hu�Գ�Ɂ)��1��&nx�o{��(a�b����1��g�#]t��7,!� n�k�N�ܝ����S9=1��S�����u0���[���2CU��f�����H�ރHb9a'.�O��mb�2�3�_��a.�lD�G���$�;��mԏ� 4���\�U��-׾��efv,(f�%<	������6����.�f��
�{�T���P!���tFCX��{�??�K~uԟ���1F��sk,�J���L�1�W"�Ŀ7�h\�#���u\��v��dL�����y���OӔV*t�Zl��|[�5ۜl�O��n���.����g���]������ŀ�FY�+9��@<�xO-a��_@�(C��:?Ow\��n�ު���F����,o*A#kFt��>G��� � \Ryvi��q���(���T���.��J���0�6{����V��M���J�[�g�"ԗ���SSAߏ<lj�ެ�S�=��8�H"�G�J٭��/�̒V��&쉡�mM��rr�T���r}�~�J��f��l�s�{���6��,��ysJ�[���_�/<6�#��P$p�$W�c;�Ń�f"`{�ج�n���<���$�[��@œQ�i���Оj�u��W���<6���4�E��u(�-8>AG�a�.G�e��H����JW�~p�*��&�㌓-������b�Rkf����s|�ڜSjQ�����~^�l;��#
*�J�;�t��~�[ϼ�����N�\�hf�gwU�S�z�诲q�##yu�b��-Ɩ�r�3��i��������0��PO���?\����ɗ��IE%%i����o14j�H�QG��߸J$U=��CZ��(���ȫ-^q�.#�<xz%�2���E��d�������?��w����NN�R�+q"���
��T��/9����ԑK�g֫�}^��G���hE޽y7#�}�8e8ߘwUH4T�aSL�ý-��Srۤ���O�^�)٬��d�E���i/�,إ�':����Y�rߩ�^�B1'�֫�Bx)+��Φ�}�f����E����
�	�x����X"5!N�M�_lv�ށ����P �A%�fL�f�ѝ�A��=*CQh�M�
E�O�\����B.v��΁�t�D\�v��0:��5���dPZ�Wu�)\5�#�� ��X��Vk�`L�J�S��>�^,g�U_R�̞͂�aIs{B����dތ�v�Y�%8^<��kb�v�9M���0b�ndDk����@��+8( ��������,�X��.�y�8 /b_3iU5U����@m���0�Y��V��E�Pm����@Ԅ[9B7.Rvj6zsUYޠ�vH�4M+5�um-o�����݋r6z��Q� �C��dq2����f���������_�� yHm�q���O�ҏs���7%�ot��}�q�7��S)2�}�@��{�2Ќ�:�R�̈v��E���b`�Q�yMŻ7�:Lh�Xϒ��N6I�X/|+d7 ��_�踗��ZH?�ޖ�D�ܓ�7���_R�������h��a��F}瞿"F�2X<7yU�9J��iޮ�%
��y��Y�/`�6t��I���5�q�	�]��nM�"��Wu)�� �a���G���Z���?wt�f0�ͻ3�E���%�P�R�w���G;_�����	���yv�	�̇S�~�_��BA����⥈b:�sC`z�
dbG�,y&;�F�%��M��)���HEK�Q;SҹU�X���8l_4n��th�Q0��z��q��(HRq��-�{T�p��jx�țQ��f��\o!dINq����!e��**��ϓo�ǉK^؂�i��j�����x_jK�V�Hٗ�k�����k��#��7=�������m|�x(_$����뿱�퀗/q�q�<�>��_뫄���|��;�&-����6���`cs�"��/T�
����￰�`��-�؅��/?�S�O��\�M09���ک�]���;�m�����2�`�2�Mek�;c�7��i� �F%p+�"��ӛAl�*(�4��?sV����c�M1����+��k�Șo�,g0������o`PL����q�6���	5��7rt	=G��c���.�,��_�������Z���
5��r��P��5��q�=�>#�0X��o>�'��v�Ծ8� �BZ�i*_� z�!tBɖQ�S�)ͦ@!�����&a�բ�Vx!�6IYR�Z����p�W��w(�*}	\<Wxn�@� ~>^��)��/�@�emX���$mg��pf��ʠP�W��5`��k�������{j��C:��Aj�tݝڟ1;颔0����{3<	݌I��Ji�}~ܵ�Ɍ'��M�O����R�u]
�����/���[ c)�%P$���Q�`I�� p_�]=!�A9�~vr�.=��hFj��Yc�C��g)�ydʔ�m��>���]�L����C���HNF��0^?B>�9mCڇ������?���ڧ�d����Q�i�˯.���C�yiJ080ArH�����5䏘-H��c��誺��-�^���n���.y3SH�|ڴ�%�WL(9��W�}�پ
���gi|Q��*��%���ֆ������{˶R]�vHMr��MΤ��[B6#�O� �t��9�K�~Nuu=,S$�V�|��}�y���0�nY�ؖzl���?�o�O���b���cG��5:C��}B��Y���.*�27_��}L圉��4��~S���zV�cP7��^t��~�\��{�̆��*�e�o'?������0k3{��X#o�0�c�����U�t��єO��a`^:�D��B��&�.��l2�oL����p�U���b+���qa�"��?�������u�g�#��R�Bz��aK~gS���1��-�)�(�9�`<3�o��f����q}�V8Pl�포d������^����uB/w�ɉ/���۬��7��e���������c^��^�T�p7J/g�o#<��@���ҍY-�μ��E0��)�!�76���"�n�锬�a�2�����ؑ軥?7���^~������O�5i����@ADd����G;VXN
�e�{�J�P;�.3��7���aj6Xsϵly׆��[�.�S����~q��������߼�>���<�o�.D:Q �p$�շFz�K���|�LN��� 4�T���u�f�e?)CkdF�a�G%B��ȭ�����#T��en{����������:�ڦ��c����B�Zk���Xsvl�Ŷ7}JW�=t�M��f�/� D�KR���M�]�S���y73އ�Ն��C�^ S#>6�'�Z���p�n���%:"�˒��� ��٦l�U�ӨP
��C�~}�} /]\�fp ��tUp��x����u[N�=��N�y�0�#�U��7�G�ܔ�o�b�-�h��F�����~��H3]�k�ڢ���x{}�S���b�ڵ���c!��{C���}@`{2u��fWi<	F3���e��x{����W{�d���A�xc(-&� !��V����X����S5qIDf]�{Jbc�������I9SLK��&���1�(!��<�TUkS]�A��
l^�+��Q������_�o��F��>si�t���) ťW��1�Z%����ã�9�z���Z�E�>]���nC�
�i��$�L�y�<����A0�&78�l�@�"�A we?�ϳ7`�K`7�^���,��
궞U��b�Q\�* ���ꦷ�V�@/ '�:��
]������m�_Qiq䖶�~��	oβ����
��Tr��B���<a<�{l��`d�YcZ���_�_V��,Ci1���x�`.���%�L�Q��L����z�k�H�x��5X��g0~}UI�qҧ�$+�D���[�Tx���3��j.2�C�r�I4r~X$e9��h��(N�ʹ���
O�Knu�jc������T�r��S�0�`���:I��9N����=Ĳe�q�pk�`	�I��2pSz���SI0�́�X��zA
@�
-��?볜�Ӎ��7����|�c���5쌉z�^��C�Q'�h-���Y,x�g`�Xk�B��
w�`�A�{V�R^K�fJ��:�K�#��� .�[��鿖9����K��,�mSfq^��ަw�v]5�mr'.Rt��U=0�K��V���s	�3�B�Df@��u���fQƺ\������s�:{`����n��G~Px�Pv�W��=���:�a~]ݞ(�3^f�f���>}��w�w�ǔ{�
��49�1Kw��xѭ�r���D�]xWD��A5�|Nj�;<�^l���P\�LprJ�Y��-����ԈS-@s��(��;�������� A������3�SJv#��A�!D+}�#6�9Q���n��?��T1��<�cOd	�p�^=::�$D��{W��ފ�-�Nq�J%��Ԣ�i��nB�H�05�U8������Y�zѽL�X�R�Mf�;�s����:������Y[4�	���w�Q�g����ʉ�6���\�>+A�5���vե�/�ɵD$�{"W����}��.�xR�7I҈�n�Kq��J�����3�ѽUYF���%���&�����,R.�����n2�C�$�9��� ��3VOO1��R-x���Z��LaC R��_�s�T�p���}�YL�я'A��V�RB��BO	ˬ��,��^(IV㻟>mCs�BK<K/B���[��z<��Zv�{���'>��""��`�����@�q�~N���Ov�=v��a�wC-�R�\�^��e�ޠ㑹�M8d������`���B��%�U�%9��j�)���i���;K�E�1SH��_�9�+ ����6���Ġ�v�h�����ڲ����\C��F��r�Ί$5����<v4����=�}�;
��{>��G.en�Xؓ%� ����\R6Z�]����K잹o��' �	�no��C���Hb���`��9�1�vv����fiS��Y�>%3f�۲�/�HdO��Q�3<�������:����[Fi�ⱊ)���u� �:`vLL.ͅ��~@����T[��`%+]��J�(�[y����%?�P4��c�8l8sj���Y��g`Cl|�d���
4��Z��Wf}��;X�.�0u<����A�b�����Vپ����]_	+!M)Ү����;�=��!pr��!����O���i�6m�d)`���Ϻ��ө���y����*�D;-΂�}�];Y1Nm?��a�V�*]Tg5��Ҝ~���+4|},��H%�j�7�!�/:D!=M5w���+s
3��A�^��Z��	�����$��̀�����',�u!>��L������24��������H�,4�v�Y�"ϊa�����S;x�[[�DյTߦ���{:��,l�5Vz�����h�L�u(Ow2ʪ@�1��	��e+#n�bL����`-o�;��%��t+-��R�啭P�+$���`Zǣ���?�Y��2H�0��]� <菥��7�p�Q���][ã�
�sBFv�	ڱe9XI��5��V�J�G�T���&�o�A���ۮ���Y{�
��ȫ����s�G�P����J�n��L��{��؍�HB"���\��ez�Y�o��p#0KU=1�zr��0�` ���k�Q���K�鲋�)�>�%)�f�A>�-i�͒:BUXEz��Ҩ��6OёՁ��6}�=�E��C��;�?�6�Ri�<i���An��z��#zQ���2�=�g�Q����]x%�n}�}��S<G�S`���(���t܈I�� �0uc�YWMoT�X_r�Ğ#���S���˾��������$����]�4|�\�������7Q�$a>d�ӟ����O�M�������H�+療����9�����~/������E�����v�����QԀ!@�3)�l����M�hw�Ҽ��Aa�<kv=:�_�NL�@yh�Tk�L)���
u4��<��1������D��n�^�6kC���wt�l��F�S�8}+���l�qzΟd�Y��t�O��N���\>�i��Lq����/��+Ur^�k���K18t�t0���p
��<���xe�a&>�"�RͶ�7�$�9�]Ԇ�L�6� �yҥ�9�o��,�K��I��-B����>��_��â�,�8�Pvƶ�����Ѭ���X�8�n�H�Ԡb�d�=A�N횔/������-%Zǁ��N��5���Cm�ĿNY�KrH�&�h5͞��f���"���@�D�������G� �����C[?�9�Zf�wXp3x��ހ��/���o��_�8k�xT�$�(�)!���z&Ӂ]�3qNL������dM%��ɂǧ�8L@e�1f ��ͭ��%;x��p�iY�Uw����+�`Wa 	���&��fב�Ԛ�Pd߀��Y�b�^�Î��z�K�8}�$�\ý���Rxy��i��O����b���������鶚����
��K�p�Vox�����.Kr�ڑwy"�Y*��(�x��&�������#�n��>~�7��m��Jn��=o�Ǩ�͆6-�2b5�;���>��?8�vH�&v��X������!�gu�I�����#t"�*�R���礀(t�c]�5�>4������q�`T�U�"�br/��w�ˀC�̝��SN+jo`�Tz�ٱ�ₜ���<��$G\�t�\As&H��4Ă��#S�tl�SI��!���e��Av窰=�В�c��:9Ӏ�[���X��AV(㮩K
�I�&vĽ6���������0���ϖF�5hd����i[aALY�b`P���0�$�l�(����Y���E@����e�E�m
�L@�悒p�� |V60���^TXoU�U�S���7��}uV���F�]J�u���z���!hr�i���d��,�cny^�t���WJ �Gv�u�ܾ��<ʚMp�ٲ��V=t(��UGﴲ�0���߇T�`�1f#:*�t���L����_c��^���L0���O�C����Q��%q#s�a��!�ʥ�#�n�E����m᪒�%`�lu�R��{��<+���U(E�h2
�����;SMcg=i�w���~��&7�@�͔�p%fN������'�}е�nѐ�B�:��G�t3� S�C��lrƹ퇳~_Q����v�[D���}a��Z*�{�Lj!x���'�6���K���w	�3"[W�h��;� 3E���[���;E� �e�X���;G2�`¶��XJ���<b]z�O��T�`����_���J/��3喯�gQ�%�-1!�oN|`4/"�VC	W��j�JÅ2��ѡ�X�1�+��*����^�t6�x���S�MFG�%�DBw�~g��<YTt����]��i�њjt�K�N�9G�υ�_���+��ש�4�ǂ�+>�t��U���%c;��,����6�cx�+�ũ�\5A��lQ�,��nF���q�YQ�gv�v�.�$�����F��@�
v1D�ׁغ�^Ch�)W	&�=�K��k2Y{���~�%��R�"��A�ۅ��^Wj��F�Ǫ�$̒!^�u����'$���T/���V�}�����G��i��"�4�]�<߂�#t W�R�C�R�cl6y<�1[��>_��#¿�_�Mf�G/+�oM�����؄�(����
J՗�72	Q%���Jo�rԼoE)i�Po�9g��b�FMs�Ø�H�����v�,��m���<�w#U�V-E	.�;H�pp�G���XE��|x�D���ǃ�x1��ҿ\�:x/E�z����d�m�'�/��BK𞿬�ै��Su|.�V֧s���'X�|J^ q��j��h����a+�����4�4�� ���չ�&�ܿ	�5��5�~�E/~k�)��o��i3Y8\s!"�ě�����B�_Zl�Ek�[u�ٺ�����uD\�DP�]�Fr5иӆ#�npAO�7
�ĽM��:b%��)-B�>��\#�Ϻ��0t�(��/�^2�MkćK�s�e�x�I|aI�>��{b �i0�� �\9��&��n��x�V8�,M�B�Q�4T
uoYiݭ�Ǯ�����$f�n(I7k2~��t���.�
�R�Z�x�<@���4M���q#.��E�R���BI��B;�a�l�������٩����]��jCo�mщ�_M��Q �Y��c{L�����-���~��~Z�\_�gh�r�4��&bKT.��-=E/��6�&s�M]P�h�8^�	���'˥D��<� $���T�Ӎ�$I���uf�v,�k�b<�%�����)$E|ҹv�9YNelS�C��Ͼ�~l!��qo��G���E�w!��3uj��r��� �g����xi��ni}��8y�N���9s���Xs�x9�boMs�Z��$E��7"�d�-��^�2�����Z}�Lĥ(��*��U8�T.�Y�S8�OO����ޥP�{�GtX�9� �$�,1o�a��l>�[)e�����4���D������H6Y�Հ LE]�xR���a��w]�+K<�PMg���'P׻���<��σ�`���]5�e�1�U�R��y�?��&d3�%�YG}+)��r�����	 TP���9���_���{��Ƥ���5&�}�������VR��bX.?LQF/��>��9Q�r�E
��mE�T!{_���T,=��<KȾ�����8C�S���E�*E���j޽�[Q]��AlYIu�F4���:�;��!F��W�c�*�
+��Y�IyVX�Pn��-�
 �A U5��oS3fe��wч/%��"T1
�:~f]Me�����If�|Q�$y�6*`�m�U��p8���t�G�r����0�����|�+b C��<>���m�{�'Y����Bd�Ѭ����T��$`�Y�e��\�'���N��]��c�FdzS-���6�2�2�:��^�PQ��Vb��9��&z7�$�`�M�f�H�ZA:*�fZ� "�g��c�ƌ
�| �Ma����4x�@�N业��6���K#=�,8[���UA~�<dyM0�h���mr�D��|��oQ�t�N��#�E[�����N�]��}��{���y�i�#�t(�Utd��x�,���f�qo����r����<9z1��-�`K$��h5R=��O@Gb ��qx62�V�l+����:0��Au
���[8L��W�����(��mH��@���ʒ-�u�oT�q˄��M�� ��r�$(���Qy��R�O�#!���𞥖��Y�\nW̼�:���=��7�t���9U(��S�бDD_:Qs'$���	�h���y�s����1�.t��&w_Jmڼ�7��/�Q��47\ �;!�Ϗ|����ڦ���䭱¦%kg��7s Q�W.��m��z�Ly��`��֐h�1˭Z���i�����5��]�{
6��[,Ye�,�J�\�@�`�mS%��[4=����8n/��ڸw��W��q�b���W������� ��f��b������Mڼ�IQ%<�J�t8� у7r�^	n\�E^`��_T��^��ʼ�LA#LF�v��4ڒ��H���6��l%e�<��s��Р��z��0�,oٹB*���[����_K!���+Ը�w*�j��J�6�6��ۈsd���`
�Nh�,�N����v�Oy/ �w~_��*�vU�<7(�Ǒm�b!S&Z��f���:Ժh�FR�1Q����)�1��Ѭ�0=�(���E(}@$'7��Y~�똊ov�$���׳�M5�o�׺��_���>�<��8��X��b��Dw�"��,sW-K�T��C$�l�d�if�Q�n���'<�>��T�p J4O*�;��}����1/�2W���䷕8p���O�Ǡ�+���`(rp�����A��K�Dh�ZI�Ӏ�.V܋�٦�Ү��8uc�%���=6h�����\�k-P�͎��4Ɯ�$�D���B#��R����ۓ���l��OyК��,@ZM���jP	�ԗ��Ͽ{r�J�y�yC��v�l���f3u�-?��!vQ$��5���cS8�|�(�-�7pp���O�,b����� ��:��2�p�A_�v���fi�XM8s�7�_f�Чo�A(�{�G�T�҈�%�N1�f�O���3�
(�ϼGu�RI/����D�#+W�7|���u���'���I��C�&wQ1}��5H8����/���s9��qc�V���q��kSP�H!o�Vb��A�tw�3���<?w��8Z7��-؜��E� B�"��������[R�e��п���w��n<�@pl��L��]V�ZeI��)�7���s��ps���0�dp��$�ɫ̠��μ����TMa�y�hF�E�w��h���,�>v�����!7G��!�Q���eF���c�q�Ƞ���X*�DW�j�Z�\QV5���0�U��!���N\�PD �J1�j!�.���>N���ѯ<u�z���t`(񛸨@�5=Th�"�ـ��܁��.	B��ַ�#iZ�����ŭ��='�R[Kꪜ2�سc2��z1��Ơ�HC�jl��L��>n�gu�qy8bm�z� ���{��bW���хnuoW��{�Ӑ������O��[��ik���:�,�Q.o��[;���=��	C|m2k��s�;�;2/���K��Q�"8���+G���@F�`<��)�3)
��k�죌آ�ƏȀܟk�]��Bh�P*
�Or	C�k��Z����3�^��A Tg ���\]p�X�~� _G|������K;Q���g;�?��oX���SǮ�u�ӟ���߇7�$�g�����R��{s=�e���E���a���w*u%ިW�J��1�5}a|)�}�aTԛt#V�+�|0e�'�k��b�0Gn@v����H�p��ܵrwg�&�8�S���"ph�FɍN�v�r5�J��#��I ��(��7��Wn+�6,�ܙk���u�=��?sph��rRfL�iJ$�^��#g�7��:�i"��W�%}O �t]�^/wj�KDh<����u4b
]m�5�<�� ƾxu�:fΧ��d��;�B�j:�� A�"��<�TQ�R����Y��<>��zl�ݠ�4G��!��+Ư[��Ln%vȢ�� Q��橽�l��;�S@���;:��W�`��t]�*��P�m]e��i��ޥ�x��E�O^R��Q�c�*yA�Fq�P3�^�%��
�;\��U'󔇂P�&.e)�>�߸[�͹��q��eV�Fm;��F-�g:Bt�o��g�fˊ.CJ'�U��[%9̖����ݪ�ԜoQ䋅��~p[�A1� �o ��a�OF�M�F���|z�/�$�yē�ӎ(�5M�"&Qŵ��9�Ho�*���+o�� ��i]��������j��ߤ�o�e�UX�������fb��dc�͠_|�6G2B�ʑ��Ay��Si�>zr
_-�|h�)��-�X��ơ����-�m#�w�֝���%��o`Ƣx�����*��'��܅h0��-f�a*k.�b�Ƶ��a�Y~/��^�Q��﹔\.���<���|���?4��-���3	f�Q*�Q������]�e��K
������C��z�-�Kj�5��	Yٵ4�nbs�]2����r|��k���M"��6V���-4f��QnZC#
��f�M�x�9��/ ��O��q�ƙ�/��c��;����<( 5
����1�Jz1�y�Qd�ݩQ��@�q����e meR$IŦ�h�˭�b�كhc��S3<E��ؒ�FH����ɚ�̍�sa.���SJ�KK#atnW׺V�E�"|*�U2iV�䏻%0�3�E����W�y��*^�Ֆe��6�e�9�%^�D��7��﯍���P����/��_��8_��>�PX-��'GMSW�<g���n�_�Qҏ���З�#�?�0�=���0,:�c��^��m�)�R��T�3��P���IR/��}��T��i�T�!k� U�,	�{W1� Ϊ1���Ioh������
����P �B�򋷦�{���=N?�ۺD
����J5zLe]~D��V�K�W�K1��y�^���!YL�z2�k@���x��UR�^Qf2YJ�ع�S�bB(.�э��ze����=v���qb�R�zA�a��:��.e��Ox���ԺK(��+�g�ꏱ�8��=�c?z��p���(~��}`�T&�<E�{>젮��4������=����� �ٰ��?�p��j�/z�!@D}�@Q��sTB)�B�m�}
<���9�O�\�����s�4��Q^l|��72Da����U�����>B�����V"�՜.�d��n�B��v��ɣ���o��Ȩ��A�8�ծ'Ø0�lSû���V��n>B�v�#cb]�LԆ�H���e��8}T�)us+�=�n�ګ�<;��i�r��8O�4th�>K�����~���۵�`?�w���쐖�OsQ�	7��Le������!�|�k�|����gms���d:�8Y�~�wC[���Ҷ�s6�'U�[�U�e���MZ<����]��X��$�4�S����%&�Gpb��߈p�o�q(o��+,�]��|6���]D��pc�%2Pt�k!�q�
l��g�<��ֆ�W\��/b�ѭ�]��hwQG#<4��R�]�)Ӧ�.6<�����K��F�����BD�叶�d�8�xXP."C�(�B͵�3u۴����B^C��:yuj+p��K|�7�8�� ���WJ�6���5�V��Aٝ�;�B����0�G��H�?��bW[M��Y��79�	M�6é�5��k��.��C�.�te<�`�������x-l���gV{���㻐�4M��a�-1C�Y����垯L�ب��o�j�����)��v%GX���@yN�k�b�9�_��Um�"��)�Q��J^�֟���>�%�>R�+� �+�z�^��T<�9�����_cN�<�Rg�P[��Ԙ�*'u�M�<����v����ʺ��!��O��i��z���^�i���9G(�痀(�����wDa@�Nd���7���u�a6%9ew
:.�3T.��� y\� :h8i;��q@_˃v'̌�3���8���A����5*�U���+��x�uޘg�u�ٳ���*Pq�%��凪�������`��)�ͨ|n�U ���ߕd�A�Y��Zfv���P�n��~9���[�P3L�2��3ĸE�;ј�
#p�,�DZW;(����F3q e���{�9�|w^���kF��{Ѽ�H[ʟ{�ߘ�3OE��l�<?�o�A��۔	�U����>��E���t�Ӽgs����!Q��~�.-�7]�c�'t`����աp�b'-����,��EJ��3�K�wjQ��w��!�S�ŨL>n���ԙ|֐������S`a)<$��l��i��I&��!K����?�2뻗�����?��d���K�}-���c�gr�����َ��CL��ZX]��� M ͥ����̩X��m0�F���6;I� �	b
79(�?��Ѻ�&�'p{Z@P	DnX�y��fR'�tJ����򽟞 �z~5��O���ki�,b�<�n���B���,&��l�J�G_�)��9EP�ă�'8.I>��b�<�|ERSa)�5V�F�v�H���O�������/��:�XV��h�cl�h�l���=Ś�_��Igqq)���i&4�47�H*A
�V�-�Ce�`�Q�$a���J�;>B����B�C�`��;�	�9��v(��O�f���5�A��#B�
���h>��_���2�`� �ER|�m���,�F��z���\��� ����$�
�iNYa�P��d?:uw=v�&�.�����B�N��8�Wz7����i3^��V��㹬�pM�*(ցT�n�����82H�69[c�Z}�`���/KYG��^S�/�tnI�&:�lRí�� �vE�R����B�S7_7e&�X�U��6WjFO�rH���j��]�U�4ka��`�J��fw�������c����!8�{� �1����3�����TK�D�T�����W�k��W�\Y�.lV%��t��/�s��d�C<2�Q���{�`	eC#@̷+�^x�h�萯����	ʡ����V���8�����B(Y5����$�on #+�u�R�</5{��	R��cX����6Me��8Ò��m� t3`���Dؠi�xl��:���8Keq�;�XL{lS[?���jn��{-S�?"���� YR�)��%:��w�ل�'�RF�8ݔ~���(�+��@��zZFl&��\_I���r���a����n�����K���=��SJ-th���(����-��L:�+)=��vŸba��������Ϻ�Ճ�n�_C�k� �׹�:s�sF`9�k�A�m1����E'���oO��(zf�4��J��:���V�ʼ%��%Zϋ
Bun�`�M�5�4ʝyT`�׆���S�	�k!z�
�De�[/�o�A�_��|*����-���<˙���5�~P\�9�[�A��&�Mzr%kM5���s��ȶy�ѴwW4�s���_��H*/db~��߆toxH����S'3^AZ��:��{&� ��2L����K~<1h����pwJ<�}��[4�G��9y����W�Q|��|��p��D��5R�ݙ��V���I�5gbJj�+���\����m�M7�������KiU�qW�f����r�䯾���X���rL��W�~�A���c���`���>�Z���-,�/!N!��I���_��M���uf[������Og|�o3m.�Ż�< ���pWԅ��������g��e�FExw#f���J��ꀎ-���5�@�5��;&�\ȧ��DT5�6���#�צ����^����hlM�	���3��?*/���B��_J��>C
i��7�@ը�;m��x�z�����i���1���r޷��|/�M�����ן�Z�����[�e�8�����n�|E5���a�9�bٴ�>�=�j�|�{�)1O��o����uk�w��߁��@���ƈJ��]6�IQ�ǜZ�ԩ�vDۉ�:��.
��&_t���@��
��Y��-qE5�i,ZLD����8r҈G,����o�	^���m����;��Ry*e����hѷm���v0��%��o����:��b�Hn�^Y���o���RI���7<���9I��z���tW� K�9��(�$w��?qP�m\�h��'y�ܻ�� !�;#o�.����W�'}��OhU��`!�v�Ԇ�^��5WfLCokUf'Xro�9�@6�Y��K���`���g�vj[�g������U� $<��}n�MJ^�و���h;j���-���F�lFO�#�/LS"��m�e�m>����rN��J@:����'��"�}�s)L���������duNz��Ǔ�����ѫ��7%�����!�K�"*��E���Q��I�w��~1T�u���AyƎZ�Q������#�G���� ő 6@��
WN�Y}O�7��Kmt��	9���9���,c�"�sn��υ�*�;T����59#Hfm&nlL�!FȤ�r�E�b����\ٝ�c�tm�kX6�^�2ѿ��J�L��/�����m�>h��V�f~ <pu�k��H��<��f���(��W���f}]㰕�V��v�8Hsb�:���ݦ���U�j:��)��Y���frN� R�hBc���3��T~{�F�����lx0ך��L!��X_���i��:q�d��IN��*)�`�����?�sr��@{
ҏ��"!c$���u�����q;~в���m.�w����,�J�8c�z���<��(Z6S@љ�����}�����ET(��)�}>	fVO��i#W�����rj�@�J�ى�
���t�&�nM1V	`P���5�G��b��%��E�R�تr���.,�~���A��h뀎�ɞ�hIE�(���Qe����
(�{l��I��m�oE.1�E$մ��Y��T��jo-�Q(��bT%?)����)n	莟���mJ8��.�x�l �QrZ����*��4�0�D�8���+��M���8u3&�K��W!+�n�8��Ip���ٞ(����"q���w8�9���]#@'%^ R�����eX�Vt�ׄ��Z^˧�z�@�oq�+D��ʪ�6B�*�a%����
�+��C5��2�w�`I=ѷ�&���<�ٞi�̧�& 6����w]���ޤ�S���u�T��©e�Z�򚿀�f*z�	IO<��w�����DLL�[B�1&��1�d�ZO��d �T�N*i���)'�ua3)%w}ر|kwꞪwr�c��B�8��� -�!X��j"���HHL
�����3<�p���C[�[�Q�U���4�R'N�<^X?�{3 @����I�Y.��U��P`�����
M'��c/
8/�0l��e�j�0O?c�J&T:�3/����F���u8�� iꡡI�:����z���b�(�������܁CD��� ���)͆(h6��LA�vƼȀ_��dY#Da�S�Z뗡ļ��*,��D8=@��i��=�<S5u��s�t$���S���p�X5m��qW�ta�D��S�'+g�-��,�h�'ڍ�G��K�bL]�<��h?�r?�S��W�,�V����#��>.F6ώH�f ��׈y))	��;�*�6���|��f_(��4XG̘Y�Q�S�,�;Dom����w�����S�%&XG ���|�r!���X7���F�d��7��m+���|2P���1=�i�F'(s=�>�dx��n�7�"�e�R
_�6������z����O	l�
E:��OM����Z�f�dӐ95�M�n=̯��Q*�/�bL�m����6�5,,%������ |M��H�!��[�Ʌ4��rF�܇���Q�"�ѹ/��A�W\)����|�֚%,�-��W�ꤦ��i!�V�K�p^�Lic��0-0�G��'"Mr_�$�֍��x�T�̵B(�����f�ّBMo�#�Vvz��.��lO%2��O��e�6���'�1��q��-��_����y���|��t���7�+9Kg������-��"�sz�ޭt�C�ǩ�_ɑwGN��@��5ΛLGϿ\���t`���I-F噇��&��sJ����dTvd�7�����ĮM���V�BmW99��<?,���§�<��ؔNE�/fIHy;�i_4�O].���5蓅PZ�����X ��>cO���������0@	Z˯*�I�i�������4�K�g6{��Y����H� 	ՋU�>7DM�Q�`$�R�G%Ki���ve�yE��v2��B2ڣF$��I���"s�P	ˊS�!]�-Nj n�ś�5��IV�D�s���W��v �#� ]]:֩$�JEX����*+�Le��>���!6Q�d�N�Mѝ5��Hb*��A�}eGS���K[�����^dp�6��V�N&���CQ�
���^�_����@sxc_����?����#��Z�}&��N�u�89�S^d��^D|gn�OHӎ�C]Su�\�����{Ͳu��#z�Tw�j�ziz:]�c�h�֓��\��D:k�( �x�F����/f��u[1Ҏ����:����._g�z�LP�N�������it7�H�^K�_	jR�@H�Fho��Ke.-��������-m�Vx�����Mr�����-��;2�i2z;�#y,��ڃx�ᾦE��ߒI�mn�[�b��f����O��T܋����I]��S���n,eb>#Y6���p٫N��`��y*�m�*�U����*6�:�}H�K�U�����!障.I9=�l��OO��9���t%kzƘ�ti|��2�x��uF��ߓ��>N����5�[Fw	4��ޮ�&�۲�Z����Uv�<��z���%�
9�]c���1�;�$���F� u�J�Ц�;�N�0�[��w�r&�b��w,�@<z���b��9�bBU���<�$��kM�ET6�0m�����\04"��N�s}��]I,��4@�ĸxv:��Ø�G��PC������e]Ƅ"���Q,��2�A�|zVq���Ҏ/�7��Xh�B#�8w�B�^����t�>˘\[���VKG�`�߻��f�Ǌ�$ؕzm��	�a��ұ<�-M��	�?>p�s&ىr�M�K���
o�X��X�D�m>����B�^.=*q�ۃz�.�I�(%Wi�B�H�>�lU�
$�8�AOOi�N�ʧ��(��.�18Ad��u�1��KK�a.�m!_�g���O�T��7>�i��.<����aM�ÿY���7c�^�Y���6�A�;l���e�D�KJ�@�z�C��{�����Yvl�&�0�Bj�f���������m>��R�L���A�vW'�.������)��Q#��Gz}��ܡ��f!�kJ�"��1~����ue�g�z:~ǀT)���������{͔1X%���}yZ��5�7��+�P�u�h�޾?t�}�U2�mJ��Lh$^��v��`�kI�����@�H��Ҭ���!�b�$t��/�v�����j�r�D�:	',�Jk�-`۾�>e\����k�;���/ވ>�\9�����!�ȣ�q[5"H�lG�5,�� ~�L��-/�貓>�5q^u*nQ��s(��8�M�Ќ�i��k��n
��'3��UL[h��,����Z��́��7,��z�ߋ�t�����¼a�#���%2�x���
-�҂�D�,{���Lvu�נܰ[��`EX�����dz�W�:�P��}�}�MٷOƐ*�c�9T�{��b��2�B[SYYd"�x�5i���f_�s�S�$�0�Q�勾� �YI��`�5RT�_������1XH�!!���}����{k}�ghDl�>��M�h�w���d���k�"�%e�7�z��ٷ�+A?������k��Q��Ck�{�ϱ�ȻŁ��N0`Dn�����>��;�3�D+"_y�=��э6�^T]�A�V'L�?�Z}�P��)f֯fu)�4�x���0�2� �a��P��׼��ȅs�y��]���������>K@��p�����9�Vg"8�>�!"�įsj�]��p��}+ J��d��1�_���b�5��
.�r-;Q�� Oc��J����<�,�b��k��������l�.)O��ڔ�� <[��H W8u�f�Q0�ݏ��̮���8]���`4~宒�d;La ��Lٛ����q���6��I	c��M���M�u������}��,���ӥ���c���W��n���*~*Q�Z���>�d�	D��V�&)�TW�<�����5|iy�48�ʟ䟩�9+S	�	&&'
�C��o[b'�q~�W��P�m�8��W�d�ߘ���AW���i0n0tN|�G�S�}{����;��B�dfx�4xJ�"G�8p���oQ3Ek����z��U>�Ϳ������^�f�;�B�j}��~>��(� ���ۉ��E���P��w�-��x��,�(m��߄��oT"��"½�)>���H�C�.Wkcqe��v�E�v#��Ib���E��G�_�D�ZG���%�z�?1k�{H97zU�Vh����Bx?V&jos������ � |�B% �+���lզO� �.8����ѝҨT�ұ�M	a��A~��ܠN*�<��6^Bu{��Xinf=��܁���:�;�A�m��d�laR���c�g�GA��:�,K��@�+�߇����%�1"w�7Y��"�����Pގ�k��)�U]�V���I=hmCM �3�*<�6��m�j�T>ϥvQ�^�A�lW��Y��F������>W[�Y�s�ZG�5tDo �?����-=P����|:�m�� .K�����'�q�Ҁ/��	қu9����.kU�rH�i���Ɛ1Q��Bm��Q�=&�D�
�'߄Px��h�G�@S���..�4�(���,�j?��k�1-�`σ�d�*Ɵ������߈܍ƺv�kF��̻޺�@`��L�$,&� �aգ�|�<B��Yw8�tt|�JN߶��~� ����{ �j�wy�N ��N�0��h�a���KpN�ꮉ�(�OX��%�<D���_�kX���(��+���a=�y��֏�S3:�*�(����J(��:`獴�W8PK���}ܻݟ�ڤ�&T�,�S*�Ng	����*]U����yD���EvA����+l: �����ђ�Mݔ��^�'�.FXu�*�X��l:�0�)����:߈��?�g�tC6���"�w\�P�(�Gw�,��N�>�����>	��KϠ�gj�owgj^P�9�p����-k�ȯd������@���4\b�46��[k!$��	� �.1�t
��MBԭ	H��I��F�H�H�s�4��9 Ӭ���)&�������������`�S�	�*F4xK�Tg���e�{��	�I��ʊ��#>����`��j�̃�MN�z7�4�����CN�
��>�}��F�v�*VV��J[��RM4Q�
�U�d��1�}�R� /�dfuL����_��U�!���H��\ �_���:e�%_�o�.^��ׂkv�JM��$	�	����L��_6�BLv��i)G-�x!n����^`���rv�,\ɫ���&�Wg�63�A���o�Nr.�O�A	0��f�f��ϗ��ө:�s#=)W8��0	f�w2���Du
�lLb+�PN'���&���6\�0E�]�1J�?W� wol�&Ī�[Һ�����Ս@9�F��,ej�`�S�$r�snҐ�Qg5yq(B���ZB�N� D�~iN��_N������ч�e3�p$�rhA�s4H��-�o83(�����W��������H���;�>cy���4C�=��� cl�c4�|�R/���XW;���@���@�Më0��8�h��0.���a�*�����UQ���(?�V��Χ� 4(cK%�!�m���V�j�W��,��$�r��c�-+��Mo0n���ٿbyI,p�Q%�7�g2�v�n��'8N�@���$���V��D�N����@"�7S7�Ѱq��O?� ��v`�W�?����J�J^O�T��L�VDN�ViYZWտ�	W�Z�_���3RP3�^~Wo]�1�QT([ ��}��1�4>O�� �-�48`������MQ�~;p
�E�9(�!�HN�����ÿ����$��V�%d�k���:8���䜃�K��1��+�$���B5�޵��w����U}3��F�։p"��\�J^Fj�^(0�2��������w��}����0����z��#NZ��=aw_ͬ��5�w82���:�u����SRmq �'�z]EY�����Y�1ʏ���
qA5��Y��״V�m˃U���Oy�Y�����s�ǁ=v�����$��Fj����JG���'yfk��<ұ�c%%�^�,�f4i�]�$dG�w�c�xJ`T���s��0-��$��o�Ƌ#��@�5�2`����:�rA�e��F����Zn�#+��ʷ�t]�Ǟݻ��	/{h�EL$y���P�]���&�;c�贏�̨��I�C:�A1J���_��n�O��H��â��]h^j��^a�Z��m�~�$D�8
on͎�&%{�nvK�^�_(��)�� �ՠ����Y��v�kP���d�N���צ7=��R.�yd�2��t��O`�Z�BޑU!��w�%�>b}v�L!��R���j§Ty8��X���۾�6�y��u�gf}-8o?<i�����͈���)�H@�Lu��d��e�Bڞ�Tn5S}����p����xt��W�e��C�>�[����E����n��c��w��\�2@��1�id�C��D�����t���<X�����A�'�"��U>�D��~~BLҼ�0��	�
[�(W_��3�ZtH��*]+o*����zW�%f~X�#~��M�ИC��x���@�������f7�5�p�䆊^C�EmX��Hh�A&Vhc�����!����;'+ʢHU���F���P�zh�5�}v3SKy�����Q���
�fI�b�̲l;|�����n_��3�6 =A�hTP�|��؊x�;� �g��}�*T�M�1~m�Z��N��t@��b���9�������B�Y��O�9F�9)���t/�2�3��;�!��Ğ'�L�(9䷗˘���n�L"| G��­E��F�
^�J�I�����S��2_P�Ǘ�jO��K� ��댍�'X}�8�)H6�jX@��!|�,��}.L������؇s�)
�H���N�o���w�ʛ3�N�Tl�c�Ș̌�>�N�n�oN�w{��t<�xI�j'<��,M�( ��]T��F�a�v���4�$��F������:�w��	��5��K�=P�`>2D,6��H�֜�����۾c���`������;�$v�Lҳ�N$�ó���#[l6����c]�5>d����M(B����8F�9�~(`�帮DI�aMI��CԨ��j�n�8����gC?sS�����9%��"��o��)�A_��f:�Vt�oX�f����h�����<�P� ����Xe</����@�P+��C���S�2|LT�#/�?k-*̇�.��a��ˌ��+�}~n�Ԓ����;Aj�l�@�Q��o��Q���'�j�ߡ��$X�r��t��UaU�t�y��L��&�bb�qK�5����!:����r��&��6����)�w�ӽS�`F� �yU<^zSP?Ħ�:�;��X��e��I���7�>�1�U����>����j������$���^3*_��gc�{�����c�eSTљ%��dk��A�͉ ��正���6�Y�?����n@yE��J2��H����X��^~����
�Z{��֌ ������t x�.���`�9�1� )� ��(xK9X�*2�:�٨V�I�����+5R���c����Ӏ��	�99�|bD����_#�.>��D4��6k��j�kQ��e��?������3��i�F��9�C���B@9b�FD�S�u�Br�Z."6gTD}�׳X�� p��ʳ��ZLhq�\"ڔĥ);��ǃg�K�9�s��|gO��\�R�m��iĖp0���������]'�&��/�����_`���on߉�������Wk���	K�N���r��]"�m����Y�5x���6L;�h���4b��U|䔩��[�j�΍�Z�����C=&���~��aǒ���Y���u�������7������B���e�u���A��k����ܽ�5Fs�;TE�<���HO�X��K(z��t�֥9F�^3�HKRG˦��-%{�@>�2쵙�`�G��[���f)�pU~�T�H:��Y1�V=��H:V�q������勒�w	�G�&|��~�/�,�^Z�ыE���jx.$8�@��M2E���Af��� <ɣ�Iw�=B�)��w���z�,c��E�Z��W���4oJH�<�Ԍ�R��̢��T_�৐�~O��F����w<���6=���Y���qQ8UG� �L7K�D"�]P3���c�َ�m���)�����C�{~4��Ϊ�H�Y�c�e�yh`�7&Z\��*�펉�������Ps]�%�������_t�F��t�h���\��> ��"� �-����T.TE$jj]QP3a�TK�/���M��- 5
�+]np̜�"���qwtTbJlN�9�=���_��)�#�L�p�<h���x7i�g�i��B@5�we���[��+�&)�{YPҪ$�z�Ð�;	��=~��Ѳ�rV��#ى('�����!�*�����O�lM��f��1��1��6�^#��>�p��Ymg����A[�L���	��UN�|�xR���{��p y�'����F��ZSwң]�
+���j;��x[\U͉� u��c���
����P9D�4­�!H�L	ޕ��AһvڃT���A�u����tK@����T�h{=8�Q/��HH[��CC8�\'yטߵ@�?`�c݄��^<�Y�QVoh9�`���s�2�k���l���>�����/ �%���ľ�M_&%Y�[H�t~�;�5��~��������H��#3T [�!�V�Yuǣ���T_,u�[�\�c<���i�#�Ikc��|�(��z�)�p2���D��L��~(�G���g�7���Gl���q'����5|�!ٸT�g膇�ꑧ����K���[4���릅���O/�%Q����L�d��_1���G�\T�I��u�n˂k��l�]vS��nƈ�u|��.`��ϊ�
x��u�-�`O��ۧ,�s�"�f�L�_�^���B쌢�K
�é8���7�W-���>�z&�Ͱ��8�Ϣi�D��HPcl#V��Xp(6d|�4��[�+e�}egK������H+hm� �R�{�B�ӑ��UAEhsk�:����bA��WwU��N"m�ס����c^�F!!"�Gd��Q(H��-��`�ۇ�a$�nÍ�4��ӎ^�g�υ1�D:��?�N���jj�$?���7Ӣ�/�*�����I�Ѡ2ܖ�j����?m���(���+VUޗ�?����*��� ;R�,$��Z�"&j9w��#&U�[�*�K�͇����c��PO|E�Xc�ƺ��.�����>��O+���b���͈K>[mc��4�5��So�M�wA�h���6U��T�(]U��:���P���Z�.�xˋ��?D?�x �����HL�VO�~ª���fS>k�[�-����p�1Xh���c��{��mV�@~�y����#���S�ЃQ��	]�������_�*���U��Ԡ)`l�(�v��)�z6�9��#a3 �6���\��N�V����G�Z~W���� : ����A�n�>������
��B�0��F\�&�9��/ankM`��)���-��A�G9
@��!f��F �풥V�Lpu�us�����? ��<�����/��_����^G 9�� y�	@F�}�=51&J�o�`�3%���Y�Il3A���I8��.d��� ���E#����9�s����PK��Ͻ�=u"���/a��#Q�3�;/qv�wS�6x\d�'W���昅��r�Y��}�}���%/U
�-LO+�09ح��dT�V��Y�<j�3ƚ��lŉ�2��(�s�	����_&Ķ�Aj�+�U�@��)4R�ϰ���J-J0eo�l�-�Xq\�B�Ht����&H��������hZ���dv�-�o%ʏ�~����H������0�Z����u���-��[��1#m�߱x�dg>��hm�۶�M-���f]�k��*���m�,d����Zb�w��}���N!ʧf�;1F<����20�8g�O�B�j�~�+1����]G�����K��no�`��56���}�!�.�'��2����M �NĞ�o
}&��|�Q�r��S�z�1T%�{�|.r��+��^'i�q���&v�<��mi�j���5"�D0RY��2N�4`��o��u�g��Q�;#��J�Łm2D�9���,��O(#��0E�G��P�Ļ�EQW��$}SWW��Q2H���&ϑr8X%U�z܅]øJ��o�>�]�վ�qޅ����O#�W@X BVEwI��\+���0�y��m֮�G-�*���mq��������Y�ʦ���3��^Û}���b_Lȗ}��gr�(��K��1��'�v�yl�aZr$�`��*?ᕨL>�c�ă�sZk�Y�q|Z��UX򮌥���Y�xd�iw+/ ���D|�dMS��v�ah��5���g��>�nU=>�0����2+)���!�剫z�m��ʧ�ݑ��X 'bX���h�])�sLW��󈣆���V���l*>~E$8��廝�� 5Z�z�z��\D���>��=L�/X��6.-�o�������xx�3�v��� �#���~��M�lG\�]!)|��{yrv� �K�b���s[����*0�!a�Jv��x�g7�W|T����ey�޺ҠB4v.�SJ{i8[��ҵ�Ţ�Р��d�ڋUO�DǪ��]��,�*���[}�mw(X���f��D?aUlD��p#K���Pv�<q^5=�$���Cc���u_B$�l��_ۢ��&Stn.�@�9�D,&6D��Wy�����(�tk,���
:Q�a+�� %k�N�Ԍ}��Uut��-��.\E�h��H���٢�!�]�a�}3����Œ,H3�礟��f�/��#(�;��p��n�!BS9b3 �k��k!��8�3����h|������!˜�.EKÒ]�C�i�P�t٤�~�.
ʱ89)NV��e���\PJu���v8H��i���
g�+QM��k���_�jQ��#G����`� 2@��B��a�Bv���@�1�V�<3�etd�[�Oin?->*A���$��HC�lg+��a\
?�Zr*�{�ks_��r��H�L\��:ʚ=�c?SyC�&El3��1�v�(�v��\��!�[�:��%,
'J�3�q+���49C%����4i�"�C��4`��a�����{�˿�:�_}MV��,N
Z��mݼ� u��������26�ѾT��eO	k���l5�h%B<daQ?
��Z���<���KYT�J ��FQ�f}�
��)&08̥x��W>���X#[�3���Qmy��E�6����]�ᱵ���?,��ԏ�n�0���$5L ��]���J��� p$M�w����Z��$pKmK�z��*XA�m�&m8sXIQ��sϦ3��P�m�;(����pVM�d�T���f9�Q�s����:6rX��X=�v;'�J]����r�ڴ��[�����+��i�����Q�����jeU
�	[�*�疥|'�򾨐EM[TfF��2r���s�3�n��dh����f�Un�ûIZ�n���2������"^3�r�rlX�y������"���V��R߂sXWV]�zwt�A��k�?Q�O�O'��UX^c�N�������-�����:���@Wu��vJ�ː�����4�T�P~��T�����(�|�eN 1؄u���_�	<f���2U�#g^-Z�����r��3��}�פ{���݌}ӹ��sљneR�־b�U����Ը� �Ą��8��1Ұ���8�ֽ�2<�۷vB�`�)3d���o�C���^~�Z�,�/���Ѫ���̯�7��c�����oJ���m�-&��<r
<"�ك$;!8��%Q�����z������1��5���~��yX��/x�y����\��Cpu�d �Q��� ڲI$e��a�d�|J��֮s�!�CV}���G�F���EVM�i���u��M�r�F���)#��k�67�Q�i��bT�g�N���Z�����y4�ݴ�ў_(���`�奓M0��-���҃i={(�Йʲ'�n-�7,����(�1ğ���&L�� �Iřob���:�{X�t�0b4#u����*?�?c�[�1�W�Վ/1,��Z�:K�%��)�B��8r��K��lz,I��{&�Mpo�F]s;�I���NF�)����`r2cl���C���E��1d�K���Ņ�)��p��̭�9�횗���SR�O�r���$�g5��5/E����%������p�x#��o��v�,�E��I�|��[̼���^cLU��\��"�3h��~g�C�hM�2��g��ﲙ#XQ��f����rT��*]�\|�e�����ോ5e0�+�O\��"wBDG�3��̪��3\O��;_�L]���;�?��JHM��.	I`ʈ)`�y����d$��i�ݷ��-
浉EUX�^�@��
�aYm&��'��)���~�G�[�=Wʥ�	H��q� �İ!i��g{d��d���jײ�0�����~���PAe5j�̷n���.d}u^�!��`"1D�r򵌍��!E�s���Ԙ�[����"��n�w�m�k�qi1��r����|�����}O���!���u����Lچ�����(뮘�ڞ�OB�P��sZs�D2G`�1��C�Nx`�S����Uv��w��
3y����ѝ��^T0�εVZ��8����f��)��u����j&ح��,w��I����@�A��]�n��<@����ʢ� ��C�V��m�����G�V��L�ޕ��7��j��[^=3jV<@rY�5����g�6�*n�m\���x:�q��f�YVaIY���RDp�:�*M���4��[:���=�+����y<':w@�l"�ԣ�Z�T˿:!7�ʨ��P�,8�{�4G���ܺ�m�ʁ��h4���A� r�� �Z��+���Y�J-�]�=J��N���C�Z&k'_M�f)�?�Q�6���CC,�帼���y�>(��r1���Z"������-n�����A��N�^Ě{I�>"q�l�����a%��J����m��Qb��P��Т����"�8Q|�	�p{�m��z��ڤ�Nj��(J���OU�C)��ԝ�%��C�;�޽�R#v�&o��3�����uR�� �m�b]h.��^i�D�,�����Fx�)���:�N���V�Oa4n�R�]R�|����7�	����h�X�UU�?Cq�˚�`#-��u=G'�Q��Κ`���r	��D��ј��hvȻ/�%�mc�(-�;�Ks�2\)3�"��av�=�g���6�!�cQ�'r����	��B���#�p������z&m�����R#�� �y����|Rzl	�o�������U��8�����fZ�~L:�?Ho�[�y86�8V�G�@����%}Cl��b��V&[R�۔/��Y�5��V���vm�8?��hR�Md}���qa��}�+[��S/��Ia��vi}�Z�� 5������ի�P��V*�G�t����^Ń��<�D�]#Y�7�
��Zߓh�^� 	�a>7;3����xN�/WHJk�/��ӭ�%ú���{�=vG�g�b��$�X�G���Fg�Y���j03�|�hS-ɧ���6E���':8�"�H�No�{RL ���=� *=���?+���c��1Y����"�G�w�3ʊ��t���除F����?/�QL���ga2,d�DG5Y[W�9W�I��|Xv-#������
wud�����Z�8�,��)�0��2�����A�����%��w�����%9 ʛd������D�5�}�"_�y�Tl.c)<Yi�{c��P�/��o��|f�}5g�nZi���p���& o�:��n��-BM�e�������H�����նǤ%
