��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��e/�L�{��1`Z�P&�f���!�?���O���2y�~!Q�U���;��@�T��3	$�	׾��:���	�_V��Q_���<	z����.���ш�zV�M6�T������~�K�d�1�������/�<�yGC��V�m�6C���J��J�irB�A�Pn�RM��I�c9���(���yrp;��������+�u��r�6A)�Z��\����v�1�]}%�EFa��������!��W�~�����B �m��`-�(�+ָ/��<�m##�T ���7لȢ�8�^��Ѡ6��dҽ�����]�K��W����D�ѩ7�3ݝ����n��9}R���j�f9��G�L��*���H��@�ƀ�x��=���qu�y��6'��mIUǔ��	��^Mc/Z_��\��Wb�(X�	�v�<�BV;ű/\o��\Z�`�z���P�׶6s�^7I��oŇ��3��<{<!�}Mr�#�E��;Gmrb���u�鬔��؊�,���L��,{�d���%Rˈ4ȷͨ�֢���M�j(y�d�틃�Q��[��b�ɶ�F�ρ�g#͛�)����c�Hƌ{�;���W��L�̡\�a�Y�B��}��ݨ��x�*�|������^BT�
V���z|lM�&k椷R%�u������]-�NJ]�-�(�}vMTg�q��`��@�w1�-C���YnB8$�ʟ�~�.�A<�
�kD6{dȃ&��0^*�ћ��;�Wb Fb����%��R����t2������~_%��I�+��^+}�%߸���w�~����&җۻ�w��?s���o�0� �Z����;��y.uz��`_���:�;�+n>�d�B�54{�cN ��yǥf�U��<�A�u`�a�>��c��2C�#Y����9�	�^,<gDu�����~´��[@�΃tu���I���D��]ok���L���J<��q�$*jGapi;��u��Tg��������?�4��ٖ�-����(;I/��L�8�(�V;����*���*���L�8DU�ӜSզ�{�7�C6�Ė�X
�
�ை�t���2%܃�,�(ѐ�:�r�
����P���0�����&��^�&�p\;"��6^�?NE���F�~+\�g>�S1�$��֯���	9�a'�X��H8&��Z��l�=�!����{���h������E����O������q@�a kA�x����'+�_sm��$�#��];��>��h���ZJ�,��W�!�P�c��tT���X�p.�� �):N�M3�  ��r�7,��t/����!�P����/ �Qo�Q��n~�`�58w�r��,f�+�ߔ�y��f
z�x翅���n	x���E޶�)��]�=��u+i?;��f��T܂b'3C�xZ����<�83�n�Y�Z0���y]�s n^�����4
y���;�nǓ��fK����V�g"&��Kȼ�bOޡ�x��\n�\Y���!�L�uV��|�w�� ��5W>V$�^i�ˋ=��%T�ɂ���\熉����`o�K�&�5�RB���T��H)�nv�=�,6ɝe�MzEW�CK����;/E��B_������o��ٸc7�p�9��@�V�X��`����k)�ښ�]�]�͝(���������Ol`�#F[Pj!���]��.h1�o�	lQ>�J�}��8R��\W�Ɍ��3E�t*s	�UM�R���v����0�������o:��n�-�����$���J^�y#�&@�m��y<��s�AI���}Uݬm���k2�iM�60)�3~,��$a`.J�|#�b���,��`�����!�;����̦��o��=����)YE�_+�w����Ёy���z+A�\��kH��T���C�5�7o*�V̋�q4*L���W���̗����9�]N��h�َ���M���Z E�I�-�'��v�.t�g`��21I=�7⩊]�ܭ=��Sf8gf�¼����	�	�)s���}o��D��6i��@4���#)��e+��j�WR�܍d�:�1d�\�u񻟌Ǚ��/ڄ���`Z�Ϳ�V�����}WH����k�E��kM��B<�	9�]���8���y�5v�9�rk��?�2�]����j��Z5��^��&�1��n���)B��b��p�&I@�-�Aw�ݫ�ǝ}w-�m2��WFr�m������_#ة]�\� ���.٪�W��8� �����$�x�t�����I�.��R	k�{��o�I��S>��r&�=��N�yzZ�_}�M�x2#!Կ{�J��F�v�}�q�_KG�w&�ݛ���w��ш� ���5��:�~x�/vH�h|.�?4:��~~��	%�06�O�~c��V��n�y]�P^S�b���-U^�u����=+�#ܭ�6J"m�1�39����<�z]6!L-N3�ZW@L�m�F�S�Z}9H�9'������6�J�U`̷o����@�Z��9O��v,)��'�'�FV���:�^��=ٜ-!|lA*������� ���ǭ.��gk������y�_6�B^P��m%��͂����kɧrDb��1�H+��Y���D��8�Ͱ<+�/پa�e�\��ݡ���0~�)�����z2P�%!R�9��A��|���[E���u>)�����P��Ð��O���"v�F�LS�h���Ѻ�c� د>U�+o'�Υ������7Oi�0��u�طZ0 �����`ٲ��2���M�Ja�9e׎���������i@�t2r�+z9�+� B�Ǡ^W�j���|�%S���sp�P�̖D���*�|�F���n���x闶���3�T�'Ow�I��Ym"Y���]�MP�[w/��7��@�G��X��+i�����-l�<�&|,c	�����D$���91�y������?i_�0&ֆ� jj��+�����B�����B,�v��uwp8��K�ܭ�Q�qf�>I'�Ƒ��4�����ε!>a�H��|���r6�qP�pJ�&wu�����"$`�(ғ4���з�:�e�Y�3AO�����]~�x~���)ߞP����A�*-���Y�cÞ��ؘ��`�X4���D�}��T:�[�	�z0;�������Q�(j��l�Ii��{�_:SD�d�D�񕡬Y޻%��'��=��<}�L���g�2�hk9P-W�;����;��X��Z�����ņ@8� ͑��F��9��t픃��eY�^˛��2)���oF��/����؄��&)h�8IP$l�ό��O
^�]/����]��J�߫r
�����a�p���DG�/5��CT����ֳ�Jj�b����m�:T���%�@@t�YrO���l�ҿ�N�>���cK�����l����Ʀ����LV2i��3ؗ���ql�j�1AU4ATؽ�[�;�����I)�
XӇ��?e.�d>>�c��m��R�eu7�i��8�v,���x��_���Ě���0ɳ�R��#	�U�j%��#y���N���B)��0��w��ղ�N��"��$�u�C!�1}¨��@��d�^�EE�N�+��LE9S�B��q������z^��8�"|t	�0	�����^4�d~$fe��_�Ņ�HZ��ᤝ��c�sj��QX�2��r��v�]���^�%�&�wH���ܖ2c�{`�"j&j��˭f}��ä�a�7`C~�Բ�옷�*�(���#+��cu1���{�R��N݃/p�g�����7<����ɶ[������ľ^�}iu8X#�:�'p�H��F��'� ��<��2L�iA~����	��[����6�R������%���%h��}�{�*ڣ����Q��4,:�z'���a�����Lݸ�^̰�`���� ��]]�Y��M��dmH�,�6G�Ä�L�D','tE�)��g�T��9u�� �s�d�Dƃ�ʆ�m8��*� 6`�f�`40�>=F8=�z2�#枏�].�e1�_��>,�0+�����<c��D�k���E�nH�^�2�B7H.��Ӎ~�
�M���eP1�z�&�GX���������
�*�&������D�e�?$���`&2�� \M���S�\�>��~��7,�Rw��{~�+�y�(��ŭСz�֥�C�}�`�y�19/���د��*8UR�C_�&efsاE�@��N{`u	C���	��c��Ҋ�)�/ԇ9١��g�~ ��"B]/+S�޷�ޒ�׳�˚���[nVG�E;<�b}��T��a��3���5�Ï����>Ú=��H^^����o��)��'�g�	����}A!��,�w='�ng<g�_+~[���Z�@���7��2���'�G<�`)��oH�0���sw�9��mΕ䞶�{�ZRqzP,�#v��$�ղ��j����h�h]��YC�߹���l�H�I0����B�텯�ݳ
b��X֚��9�����2`6W�+��i,cu2H^�Y��Y�����(���b� ?����DLB�z�NG�o�
]��x����x�*̛
1�,�-���unX��/v��ȏ����R�J�JrXp�Ut�,Kd}	X���X�?�rNg��IҚ��w�P�[ϭ٩�W��P��	D=HFs0�= �{nf /9�h��S<^,��Qz!e�G��%��4��,������<�$k����ϣE,����{Z
�CW,�'N*L!#.���Mު [Y�{&J�������o?�̾��ǢxE���18bD��E8�x��e��ڟvk�1xe��ɤ�S��ږCm��1i��ܸD�`�>�� 1̳�R�H�-��Kn��jW��bQ��R�>���7�/U��N)&�{j�������!������h/~ٟ
�3i|�]�����y����!6�cd��j�Pk�\�|�tӅ���y�>b���B8p�cwG3��ޏ�"��U������@H���CX�]y��~�����Z�V��W�FW��Yƾ�`4d�p
x����r�=�!��pE	��s) �IC�й���6����J���ۉ����^Zi��&�%c�_^�W_��|���9�^�-���|r˿��[��Z��/t���L4S?p�n��e��8gG����PV���W��\�����B���:��b�"�zvi�i���5#Gab��H>g������K�s���mL�;��������e�r�����Z#�Zw������5�_6��։���'�n�k?.���b��(��ǐ�ЪS��`�\�9w�l7�A$��*MU��f��z��ܑt��+��5�`]�RT���w-�qtO�A'w0Ap�$d�z��X��ưԑ��^�<����OA�U�#r&G>�6�RȋzK�x��I6��L���sGB�ϯ �/��>��ž�(�^�zAY�rؤ��	�m�5*��!�P��ӂqvF�`���0"5h��Z���t~�+���_��A���!��4�-X�G�E�"�386����"h�IlV�9�1�FiH��9��ծ	\�{��/k��~/���~�q)��pєV��r�����i��5��m)�1c�@#"EcvY2%:*J/+OB�b�9�`t�o�m�-f�J楏"���Ϲ#��ì�XgA��e(������'�&d���%���m�e{���%l��p�V�ƀя#��Ў�����ʤ��^��)!!�Ŀ�ʥGK�;��A��M:?�2��)Լ�WA���R�C%\8�'�^�+Ѱ��^��"ՋE����Ʃ㑸4I�����$�u뵢�����jW��O8�����o~N�d"�JzА�g�ҡ�KKZ�N\��+��##�������{��2y�ֵ��y���R
DM/��Ԇ����<�'�Q�w�G�@<�j0EV)���ș�/kj��CwyR_�Q?k�S8\Z���� ��w�Lmn�����#kqy&���x��w�5V�x/NWj�L_��R��s�#Ŋ� }/�a"�"v+���������b��������T'*h�$��ln�lKb���:����e�fͯ�����^��@�h�X�,��q�������f
� �M�3��xd"��v�����t��*,e��%I���$�b��^�-�64�l���s�v�S3�=)���!���2%�Cǉ�E��ʣ�[ l��O��� A��i���!�ùV8!��=���淝�b�
+X}����D�����>!��i�����՘��W֘j��EQ�"��-N/N� MF�/o�`]��.�\���|�5�ޏY��tXe�U�����ূA��XX�56��L�3�i���]p�ܼ\�6��v�`W�6r<��<]�jm�^O�w�_�>��f��j8No�9P��A1��o��� !ȾΝ���DH�>�x�v�v#���j����B�n`lX�|$�M|���n���)�i�Iי�l� U�;�0���`m�<bA�˫��v5o�C��v#��2��Y���e'����&��t{����r���&�؜of|�b�#���ڌ��vġ.KDGlk�p�:Q�{95a�v�}m{�Tc�^
�bh�-�I�3F�屒�d@��x���(��V�B�|s��y��x��"�̣���$���[�^����"Q��KE3��ژy���M"A���s�C`�?�%������/A� e��g��ú³�ᠬ)cYI���;cy��,�Z��;DFy����ihMI��<��/��|���ARw��P�I��Pg�JA8&P�a��
{z2>rN�=�JlL��;WԻ6)~?�qA�d�[.�Ƃ�C��K�X�i?�"c��N��BQ��Y�]��H^ RX���6�vz&��h��-�1!�W[o��g��Q=(��P��7�"!��]��y�q�@�yu�ؠ;s�Z�uw0�O�b^*�����e�[k4|�����k_���Ge��k<�m�uk�K+��J^� w2cL����`�������zD�⤖2U
�7�u�x���� ;Edjr
�mÙ��yFv���6������
 2�HP�i��(���Jq����F7�� ގ5�Y��v֋��ˢ����n��m �8��-�[��C�1�} @�'�>�IV��
m؞b���d�+�.����?}t���ٖP�$)�`������M�I���e����u��6�?{3UQ�i��BӠқ1�=�˹(����rLH�.�+(�)L�CN9>�X9��nη��i�f�%��S�w����Az^�
��չ�s���ѡ�6d�D���9�E�F]��ȪQ�"\w.s�܎a�T���<���_�5EWU�s�ܚ��J��݉y�N0��������W��o�� U={U�зu+V%W�Q�e����U���	?�Guث���D���;�=A��ϋ��� eJz@�� 5�1�~��\���c���
6]*i�Ys����:dΒ�u�_^$pupB��h|o�0��z^%���~���������g���C��n�=\�}��Ǌ.�_��!�t'��2��}�����s1��{+��"�>U�Rv�?��Lg�w�Nޫ��# ��|�|��6d��$F�v�)�� $�LX�z�.v���W4c]�=_I�.W����l4��]�ɶ��r�v� �cx���l�K�G|N0�	�I&�"��~5�<k�ά����-���@�f��l���=G O���`<���_�lh:(eص��6@������!�_D.���{�Jӵ�g2!ю�,��Rq�fD8�AF�x�_]�ЅZ-�CX�2~�.ur~���+u��@��颱�� =	'9���������>��gӞ���|���-��V����K�B ��N-q�m�Ï��-��"@#B"�!���J��8������E����ѻy8�����uJh���;��;L3_�v��2�����s�A����\����{�wq��1���+6oE���Q�����Em�";'���)MА{)�S�r"�"�'˪)G�r����сZ��$��m}�r�3�j�p���љ���"壉��y ��*��Hð�%܄ L�@�{����ظs�]��g=_�R�R��fn���~��T�A��І��^�i{/��T5W�峕,f�#���cfL��%�!H�s,nrJI�걦܉� f�m��ꉋ%����Y�ڽ��� /^.��	�gL�
Rh&Ǒ�G�La�n���:��k�\��K�+��dc��45�:&:�%5O���$��/WW	!�y�a��~��4�n �����:2Vz:���A�����7�$
ݶ0�T���_�xQ��)'o�=�I��_Z���/~xA�z�[v�s,;�߹�
��\�B����'�g9KB������O�M��V9�r��6���^����Y��a�)��9�BŴn��*�u�-��ntG�
���~��f�}Sm�$�{�%��-��7Φy�4�a�e�d��ZPgg9q��!����>�-߯��>�!f��K'?0�Ƴ�$��ڕa� o�dm?�If�2m�������t��&`�RC\=C$�����!��ݰ�u�о�ߕ9�P�\�*��9Ku,��ٯ�t�h{�d�i��Ѭj��<�����" {)�a8_䣃���^u�f͠�����d����uN��g�ظ�9��k^��&����N�Q�9���Dg�~���4]#|�D�5A��k����'����	�M�a$�j�J�m�ˎ�N�7��9�*ԑ>�2��P��۰��'v��X2~x�B`��u�B�P[n%��J�< kVA�[N�^��CKl���K-�?~�N�Yb7�E�ב�핼G���� 9hǅ�c�y;���d'��%�b��9�V��&�J�~����n�� ���z�6Nt}6��O|����ܛ�|>�Z���[Fa�{��0e��\V�=��Z��>�T�{��鎊�t��P9d� ��aS����)77ϐ�{Ώ��d�!�ai����x�EJb#rQ=f5~�S�Ʈ'Ľ��"`�L4`~c���.7���j=,Q�Lc�Z�!"��m�/�*�H5'yQ2}�i��d�B���`5{���qB���c\Ik���n�ey���O	?���MS	��x�j(�~���"�/Bݟ��EOB�G�`8�[˾��}5W���9��i��Q�ۗw>ܸĀ�=6��&��W}�wj�t�M�E�؎P-�i��znq|2���Q�a�����5���b�lk��W��`���������RMv����"���/@����T�u��;�V��%%��׺�@��AZ����Df-*�M�XMЄi��J�d
���h�4D p�C�0~�@ɭ��1���-�}~�|�����I�>�)�R �, b)�t熌�`#g�Ȳ��;�h|:ԣ�x�f'�2ݾ��@3)Q��� �}�|���w�АNG��Q�B�� o1z�Tz�jQ.�(AD�T|���E0��u�u��k!���a�6��y�����ṕ�fՖ�:$�֜Gޚ�Y)�A�!���w�т*=��k�FD� N.��&��w���E ۬�O-( ���+�����=�ɳN�`���-�$% {���u�[��zgJ����=P[��/���q
��["�^�.��d�q�2�h��J����3Ҧ:Sn|VB���9~��-�T�=#�ŋ�'ɷ=��/�~r�@C���rV��?����W~85^��"�[�e�_�}���~Q4�Q��ra�p�]w2D��Z��Apԝ����Lrh�������Ԟ���N�eU������o�6eoʡ���f�$�ưB��ڂC��Ƌ��Ĭ-�. �?+�ɽw�7�Ϥ�Q�T6���N}��{�������'�쪹���Ũ|��䅒�983b��<"��U�#z��!z���U�m9���0����s��:gi]�ئB[�S�W���^�ާ��ۗ. +}�֨���Z{�L�p�Q:�]Fؠ��UOg�F�P�%��R1e���4��D�f�g[�k�Rߗ.��렧M���|����l8�I=�Xg�ϐ�ɴ�tf��%��ȩ������0F�W�Dr�Gn���}� ݛیU�S�Ť�ޭk�ONєK�/��9';�:�=�w_�VK}��Z�!��8����E>�J���S��%1���".5�ZC�w���9��Id��ke�-����(��PJ{���3�J�i�J�F�����<}l�A:�;�+�]�=��>_w��_Y�e ��6�������°>�����&A�7kx���T������=)�g
|��5�"/2<����1��5�B[of�@b�}��q�G���mL�k0�=��F膹A���?�+t�ϛh>���i�B,/��� sր�Olm���Gd�7}*��`�m�ͪ�ur	����<��,��l��ZܹC-���e�d,��!l�Z��:#���̟u�r��xsI�d��6~�m�q�9��k��]9.;�W��!����������TD8u#k�)�v��X��tyE��N���3���L�n�����;�÷�ܴ������_�މ���{@o"�K�f�Nj�Z	 �E��Si��|(S7Ni�t�8�Eų��n���6�FFi9�DVN���[�B�6��ߡ2��F�"�`�Dx�}���U0���r��7�Hv�&����;�X�^��ز
B�zk��8�Ϲ:�rW �e�˦~� �u���AZ.����>^y��06�&�ܖ��	!�������+m�8x��?�H����^�q.D7I�)�Oݟ5�U�f�ߕ���B�.`I�ߕ�@
�lZ/T ��[k���\<n��lc�?�H3 yGpX�����Вw��ҩ*dLy�J�cKz	�n���)��
$H�گ�S��x��{�t�(אc2�\��?�H�گ4@q�w66B��8ye�1 �	e��
��Ά������ ���� R�|��;�Ƭ���~PM{fp&e���귯��s`׫H^��D:��N�.ۙJP@�,i��n&�,���s�<7�m)*��L�a�U|���.����`��2�uy}@�U%K�v��C1kƊ�|Ʝ~�U�QZ��+px��G�2��=!G
�/٢��z�s iDI�|�lCv�}m������P����肠n*16��.�C{��6k
��>���

7���=��\A�َ��٬O��٤�U!��r��9$�����}��;��K)�d��j�� N��I !����	��@s�|P��^��`�M��`y](:�F|=�;j �QO%%s�D�Z*�~���+�my�t�����6ḅ�KV��K	g�9�o�Xy�U,E��� p�G+$ȩ4NA�*���5�S9[m'��p��rl��DH,����8z��&N��մ��
��ߧ�b\]�1p�|���m�2�@Z$���$�j^�7d��O��� �	�67��b���v���U�8hl���]|����	����|8p�P0Iu`7ݏ�=�C�BJ��cB(I(�2�y����6�<)�!���]�� Y�ı�:���h��v���D&�ɂ�Z&Q�&J�\��4U����(+���w%��~m����~`��>�挐�K�ʳ΅=�{-6eT,n�z�,/���8	|�;��RKG���:��s���]�&R����%!���2�G����3�B�%`�Z+w*�l.�P:"�D����=q�:;��Ă�Ԅ�@Ν�rj@ͼ�_����E[~UN�3d�J��g!�q��^�L����t��صd��-I_"���VB~␒ᦦD�P��i/ά=����V����w��	��_oX |�*��Ş��@� �ɖ�w�=��ilq������#��>J��/6@���۵���0�
�V�@�,���!5|w�|˜A� A�<ۏ�[l�TU"��_ebH�_R�5�c5��
���[i3�\��tf� ������{��KՒ�A��U/c�|���KF�����$�������.�=]�l�jAv@�wJ���#ךRȩ��r��?{��0Wte�r*(%yIiiz�g���+�c�{�bX�,��ގ��J���}{>q��BP������Ti�!�Һ�
5i��=�xW�s��E� �#���S���*v��y�5�φ������{+��k^#w1]6$���3$���&�����Ez2���J�.���q����Ex����W)��~��^r�Ƅ�[K(�ȟ5�;y�>d���2>`�0֑��j�v�P?��M��]����w�մ���K���֒ܦJD?�&�C~��a|TG$��Γ��:�b �;A�K
�[k�Y�-��o����G�����׷�Z��{� ^]���22�.Hd��%����k%!�&��f'���q�#Eɐ_R�B~w2���	N�X��9�tL��X��D�_y�HB4����y��{H?�!��?��ⶳ�U����u"W���9�k�Q��L�f\~�*A�nJ:��3�m��Ql�������xe�w�7rpˁ��Io<�P�[��������|�$��=fd/a[ȅW|�G�hBg�
m\W^����gWB[�w�AZ~�DK��z��� !FS�/F�D6��
��\�2ܜ�:�����ys����U��7E G# �gX���uV]�l��E$SL�4�>tt=��??�1�Ё88�;�Z]|mϓ�i(����:�)���h(2Zv	4� '���}��k��V��Vқ����-���֚=MD� Z2�b��~����iئ��f3~�.ա}cȢ�z_�,S=�3�����"���ج4�a��'޶J���Y�p9��Ҡ)AGJ�%�s��'�ڞ�A���z�x�C�������wn�a�ŕ����Q��
��P�+�¢��6�?ev(o��wJ��x`,[�}�7�Q e9�3��DQ4#�����/���ڋ_�'~��uW��Aʊ��8�����j�?�f�J�l����K�kv�l��"�-�)G+h�zф��n3���0.+/��=�����A	LH� KD���h��sZ�n����Y���%���>�3�}����B�t0����{��,�n=t5c�>>9��»�ÔR��X o���b��;.�z�G�Y�Nw\�-�[�O͵���lI׈�s��j1^N����:��n��Y�_z �M/��,��"��
=t4�(L�*�k�E�D��r��x8���$�5���Z�v�W�{ ��;�UtB�����[C�bL�K�0#�D�8ѳ�|� K�1����Tc�c{�9��s������F�	�ԝ'jʊf��yQ��6Kf���P����v��B���\�z?3���K�E��·�OR'�lUۋ<�1��>�U��X�^����^��>�f���#S �D��_Nr�u�Ԅƭ���Wv3e;;�%��y~�H/��82�\'�\[ҏʄ�-Տ���wѨ=Ot
\�85	*)8����?�R�Ҫ~,>��CU�ԏ�ǃ��i��H���@����/����?P�&(����МiR�Զ�=7J��t�[��-�=�!���<�F���5Q��Ğ�|5���
g�%��*��������߿���e`��}�&1�t�c�V��,����+�U�����*0�)��U��;���&佝����)kf���fwX+�:��n:
�/hTRRjŴg�� ������A|\\��X�@�����St��SV^7���
8���/pO��b)�`9SQ(r��A� �i�XU��q�����^������4� 1k��e�-'��2�4�^T���KO�bH���8��{P#_�(�Y�|[oR"��0@��Q���M �>{��eTF2������lk���7A4���G5u����/H>q(0>����ݔ=�ߡ޺��|=*V�f�U�B �@��tS��X��`�Z���X2�?(�C�~>��q-8���gTw�G�!����bgI�	��n�E۵ ,�����d��#!�[0�
��F>9����Q�J/��S���bL ���0Ux:�d�$0�P(F��f�<���ܘ�E-�giK%���Fv�1�$P���z��-�NAaS��m $�ޱ�J��K���-�Ur��FPZH>c������Sd�"Њ�</�AN�K��x�u,D��������I[є��'�o���oq��q�8-Q�Q{.{�]�,���э���|�Bz��'�v^g�mVu���ǞN��T�%Ym
�a$�~��<�^����UPyo�z�
��}k�`2��݃`�j�)�M�*�k[qt��˧멱�5�1B�����]rZr��ةM��u5thYe�FT(!Mh��?�����Tc�?��#�w��%�(:hGT�i�5����Ճ�!T�ߪ�aI�A���1+I���}P�fݒ�O=	ʮ��S6����v���m�d��{�Q�ȫ�=��j�=F�����7/�D=1��t�#?���o$�N�5zc����Y���q)!�q;��_��f}N�'�ی�o�$4�;nW~B��Ϩ�eql&�����-*-�{
}��G돲�#*ӻ�ކ�(:����P�`�7d�b9�	1�\�#$w����D�$r
��)�,�z~o"֬e�0���S$N���7��_�`t ���ɕ�ʃ(%���E����3&ȋO�,
�lR�����E���A1���Rf��vτV.�u*	Vm�Pt~[�̫��˨�p�J
���W�l�� b�ǟID��c�%��CjV����l+n�̥c�`�I�޸������'���-,���i1���w�9�+�@��9?���p�ɽ��dV�D���O�RdI�Yk����§��hI�S�%Gn�!�b��hu�n�U��-�dn��.w H�/�*������{�^�!��~�cՂ�8��Y�!*�a�kE�_��W=�%�A���:�a�����E�������DV��=6!�W~�.S �Vn��ˬy���_9e���2�	�����t�{)�-*����*����I�Ly�MyC��2��5}1��N&����P����B������wt��xӆ������h%t��6곈@/�[H����w~5g�����!opc��/aG8l�8���_��@�u�6�I0D������M��8�Z�W>�ۅ����-�^_�-�Pɾ��ND$Ă�g���|��J�»i5�F�*��J���ȯ^T�V�����e���ni\��fp/�	6Y������qu��7^��f �!^��[�K�.G�)�9mzvg��7���e~U�]�1e�Fț�RA�5	Ya$ɑ��*�s�2y�h�?�����Tbse��x��j�����L�©�u]	{���O�(NOO{�)��zv>��H�p�|�~�F&��W��w��D�ƹu�����ތD�p�j2ꍳl������_`��?���~\;S����m��$�&j�يF${�����P>�p�
M5m�캒�.zE�5Un}Z5���/������";��҂��5Ɲ�Ptg�*�5=-�zt3��VÆ�MQ�@i%��D®�쑎7�O�+}���������#-
o���� \_1�a��Z�
���ͩg8�K��9�QlI>�s����s��w�O?�;-�G��=4��0~�!�ƕ/'9,끧1Mⶬ���j�� n>��r��ct� OT��$�����%�l�q�C6�G�v��>v3c��p�_P���,>@;N�u�{��fp�"N�b5$4�Y���y!�X[PJ`�g��BxN�|Jf�2b=K:m!�b1B2���yt�����ۨ�S�ĕ�%r����g�" 1�= YX2��xm�:�xc?�����HI�"̈́�⹲;�,��uz�|��MI�]��y"^��:1�ޒ��;����E/b�9�=Tц($�4�E�@B�e����$#���_!t�YtC# �p"o�:����vj��"���x�*S�%̼7:��Yva%F+�U?p9�? �r��|I��k0yl��(�*���Ii���j��o�nK$��=�N=�3&fq���/9�p?Om�e��Bs�X��^�>
=���%6K��8l��|�d'�{�������@�ֆ�$t�ڈ��5�� g��ҥuh��5O!΂�Ek5�B�>��a��k	T�}+E�8t�H������GqEJ�"�!㧺��E�P�O�~�������I���t�f�cM+�Ä�λ��%�}����
�ŊA�|&�Z��Jt���h(r�� ^Ĕ~]bF��aP{��Q��7Asr%�w����b�c����GjF2�'F���$�}�{۪���S��F��S0[Q��,�<g�����v�K�Ƭ�&����1] iO~qZ��+o;Ѱ����J^���}���n������x�h�%�Ys�f�ꬿ˞�'h�_K��2�FQF�aD�$=�Z�Z��G$zи��,.텘����5�k�f2���&���ޤ�6����x��{�MdM8��8#��5��������Y�/������I]F�ޤ}3KՐ��zZ>"/�N�\�w����n*A�W���V�[��ë���'��$�r]�!�%a�j_dy.�bH�Zo���g����ߨ;��t����H/����*���]��au�jЃ�`ڷ�Gm�}��SM�0T:�+��G��j�����^��2���|z�ޘ��= ���cƺY$���L���2��.�z]�P�oP��#�|L����
�+;���S���A����ڭ�M� �D4�L�_�N�I*���*�2"хo7�l�k#-��6��ڔ�۾�h�a}�%��	�����j~ѧ��N�v�JW��Ǜ����������g��&I� ��u�9��9�"H��y@KE>�����E�n(�-�Ƚm�BG�*U�y�ě_C[�̤��B�n:�eLV����*�q1VF:?��Føc7��4D��� �@k�<G�$v߀/x�D�"��G&�	�)]�Ƕ�V
\�����dm��+p��l%��{E�l�;���`��g*���y���x��g�m�@y�X{zx�|�����1���������J�r��O۞�b��v.C����P Ԟ�$���_�K�IV�Ӵ�ҥ�Кcq��=��o�wYhn�=*Щ5Z�OM�M�9\%d��Rώ��!�׃s̑ ���獄U�O�u*�8��6}�t�{�H*uE���^j��"�M���8������Mt��ua+��XjUT�P���b@��`�
�fX���5yKU+ܣ)$�.�P��*��"r��/
 �am)����j��PK��ב�4�XZ��,���d��^@�O�U+	[q �D��Q�m���>HI�?�}N��������?	����r����|]��d��m'�ʛKP�;&���,��y�&��^s8�duOa��(�����`�[�>m�����[��k�1�n�Wi�	�f�H�؏��/�����P�$�3�������}��Ɔr\dSEmHPA
6�s�zG��Hq/�B���
���&~Xģ���}z���[�WiL�h	�jLf�ױz}Ψj��3/��̮_NHR܌��	հ���r�/����t |k@,0�C͵�u2$MLT�2?��UR+�����S��'�1X�/,0|?�9��D~��y�08uC�&ڂ��hUx�b �5Vl������k)�X��TeM��e�r$X+��K�rV?�tї�� �*�����6��FY�[wA'�I��A�k)J0�-Lh����L�s��,���+Q�?�8�2�� �xSWLZh����.>N�� 6y��0Lf�3|����ԥ�e@�+_Iq�=��@H���u��QȊ(x�|���՝|�c����UT?8���m6��Ň,�g��?M��-��ߙ�'N�\s�0�ƕx��^�C������xV'�Jע)λт�?��ذ��OH�)�FI�8��yD�[-s��\�j�k��.�:�c�3Y��\_5!�p�%�g�I�g��E��	Ƣ��E����L�^�퓰��cEHۿ��D��/5(����>J��E��g�j73��Qe1)�^6�1)�F�_/o I}v��n�G�A���!p)f��������1@>Xٚ�:��&ʙ����C%���lW7�O�����$N��:c�s�,�i �g� P#��Ò���-[4*<	��:4�mG�xٽ+@k�Pvf	��ȯa+9r$�O�]�����$#r���w��ݔ�Pr��~~՝EAR�4�Y�h�ݑ��"�����'�s�����JW'8<����cx�n�1Z�҂y�����Q����mW�u"�\S�{�2�ܘ��r��Sn���*E�f�lU����#��CF�?ICV��I-Ǿ,����7���/�&���XR��m��v�EƗ�
ʉk,0�A���;���������2ČVZhyp���|�[��ư��z.��V�c��QƠ_��&�giӜ��)�Tj�q�^Z�����]8��Я�#�6L�i�F�q9�6ǐ�]o��OE��YZ�B�%��'7���:e=�B��U�����D�ĝ���Y4"�V�n_A��\GpR�ۡ��[-}�+��gGź`�����!�g�m\��a�A��LӤ���{V"=]~�9CmD�"��NqC�L�]�ᾉ�p��+3ٳ���u�"���O]?� b	�@�8����6
;�<�GF)	TPe�6�.)=���5wd��r�Zɩ��"� BH切4v�$�(-V��G{|��E�w�	���u����B�D��I*�k�k\˖���z�1�ŉ���.
�R��,��^�<��?�����A%�ȼ7�+���F�o�����L,�[�Q,�T�Չ[��� �j�)�����c�c��`n����΀B��c�5'�\�����%��O����|�e$h��5�n�b}g3_ۣʀh�AE����&�}w��k��
SH�	rf�ܽ��Z�8�}��4����,�|�Y�o��X{tȷ��]y!�{!%�����(��բ��N�[�ۼ�ϣ��I�j�\�aM�Ӧy�y�8q𥅨_�]�ѭ*�jͷ�=����PA���$c�i;M�N�a^\g]�����l�Mʖ�l1ZC��]���rl���_��+G�Z�8(%�����@�L��7����: 5��2�$c���\��6���gY�Ov@��S�&F
۩�~]d+<�(8e�cm�}JkL�9�꒲��~XZ� ��,0n~���Z����r�>4n��X4�_�4+E#�����8���S$����t'���x~4������9p.�^l���F�?����~MiV�G�㶜y}p�w��g�S��m�R�x�V�*��-�H_��qL��c�G��e̬�_wy���Z9�R����eR�!͙>��%��/�c2��W3>�¯�G�P�:߲�������������?$�`�ܵcN�������O�7Ձ+��F�[������� &́t蜯�,9���2P����u�N�)�3k&=cf��������Dk�+�Z6Y���
���;"}l�E�j��hR|o��.6MZ�)��3G�iB��&c���R����5�D\�q�`+�%��}��y�zf�/d��&�� V����)�
 ��� \n��q�g�5"-���?M�IZ�����
�{�g��h3G�3j|��{9�
��g�4����ɯn��t�iZ�=��nl��~�Hl�1rӊGu8�C���ݹ�X{���9n�6���O�i��J9�?e�C)VѾ$�cǔ�� �+�CѮ7GP��÷��Kb�3�_ݩUi��y�`��31l�(�e'��fl՞ z1U�\������#\�uj���C��]a��o|�3��b2���W�M4�*�p�#nb\�G���/K�>.�*�}����A�+��h��و�[��7��L7�<&�jW�oh,W+7�����)�������$I��
���'��ыY`���BmX�L}�W�X�;�� 靶lDɶ]��'N�z��{�i��j2��)�ˆ�Fސ\��(k|(A�.��VK���pC:]⟔�ͬ�ۊ<8s�2�C>��7�M���p�jh_'�5�����G��Ԑ�j�M���Ө�~�]r��[���/�086�LJ�����2�c1��L�f��A�NJW��B6L6z=6��-HHΝ�)�V�H=v�*�U��(aܳ��16)G���9�%�M��y����~s�Ƨױ��3���<B�v��$6��ڙA
&��/<�8ĩ����ȴ�UH0�l.�	DFP|}#���g�I�;� ���H?�v�^i9)�@ȧ�ipI�=!݈[���Մ�qf��JU��f0ο�bk�A���Ԍ{�����M�.�-tСNj(����� �	r�����u��������Y�Ji �E]�a�Cv�V�{se����	7*W��xP�N����GA�~_}�����g����g�&�\\��|5�>����*��0�;
��"A�O���r~�?~RM�P�SїOz��"�����D���,�=� +��(�ܜ�Y�����X:�o�:����#�9��5�	�$�HR0����<i`P�fz!<��-�Z�Bq4T���*q���"�*$�8���Gj�6f� �ન�cԮЙ Ÿ�;�T�d)z���{��RB���ܵ���&C���ߏF���{x�P@��rg#���q��]��46j���sp��k.6- �g�]Y_��S�V�3��fn_�Ȕ��w\eJtu���U�k�_����M6�g�|�`�Ƚsh����#��,[�=�7�pU_���*񻹮�?��N��s)˔���� k,�M0fB��}w�Ҁ>�Dk�/w�`:��ZG#��1�eޤ���y��ՠ;.ol$��|���ւi��vXq]���_p�V�\���9���M��������k[�'��Ң����H���Ծ#7�:����l���:WmLqZ�������a���P����\��!r���g���Jg�^�;�rM'�����n �'�P�vɢw[p{�/�,,�Y���Lok3ro�=rŗ˹ݩX����>��UfU!T�����$v�%��{u7M���|K
P�F����j�3��)38����u^��^���8#�pPB��t�L Ĉ��"�����E��N�m��.Ape�#R�ظ^v�O�N�&6c��L�..��ȘC�T�O�٪�,
@
#��3��LM��~i�5=*h�`�1$�~ن��)Ϡ���Ĥ�{ՅP���p�Kh1���m�ټ�Z�g�Z�͐�
���-����ѭ��O,��M�v"YJ�`�%it��w��p��D���Et�$�)H6�Hp��G ������o���Ttp��Y���v:� �xaw��飝\7��(�[$��LN�@d�o�Ɓ�A1��b\1��	�>о��WC����Jꛯl�'p�"@��C�
�f_P�4���.q����n���N^� T�J�3D��k94���W:�ѧ`�< *!����gU�e�;�	���>L��\mE> O��I��E���3���Y�{����rJ��
W���T�W:�e���ȷ�0��DX�vk8꫑�����u9 9l������O�+�țF5f��6����sĆRme���Rڢ�qe�Iy��	*u�E��G���g7[�v��U���~���-��|����W��(�%�L뷑��
�kg]ᑏC[*��J�<������m+��K����E� ��$�������9���mw�P��g��r��&���>�_Tt3\B��$1Uɜ����o�~�J�s�LO��1���Dk b����^+J �7-�yb�Q#r��K<����"�J�R���P�PBW�0wAL�deCJ{!"w�{�������bb���<���]�E2F��B���M��|��àE����� ��-R�1"�p�6�ˇ ����#-i�pT8�V̅�-���'�LI4Z���^��=�vqD�e�s���@ ˽�	�66�S?����4��SЅ�Y"e꾯0�P������gI���1<�T
�RA^����0kn��pF�y��1�THo��X�Z��=�_��I%3I
j:}չ������S'�������<���i���1	�=d���ݨҸ��s�6Ǧ�������<��I7�j��\wYv<�؇��y�h⠀���O}�T����1��}��ϔr�%���(4�\e	��Ҥ�`Q�_�`�kxga}'��ѝg(H����Nn��ɢ�)
7T����41.BݱDE�%�����KwF�f�Gf�8�1�`��Gg*��?�v=dc�N_g�hO�Ž�'Z���V�HlB���)_&x�;#�h��4_����-�b-�r�w����=�f�>t]���c"S�yg�̐�[�D "���]EȀ
$�E��#�	�w�@u���$�j%uj3^��xev�5}B+��FsG�E�r�0���۱��5}���-`rC�6;�5��� �OK�����~��H"��i8�\�g��!��̯�S��:`c��e�љk��2�_8,gH	n��¯A�ˮ�z�y�t0i��N�	�70�F�l|(-^t��Չ����5�Ṽ��q=^}��~���f��B�-��7U�eK��E�B�z!S�����P����&�&ժn���y
J�p�"�xXP�.?���=�Hx�Bμ��>�P�<�f����r���
o�oJ�k�f�J˹�p�<��}l/`|�ԌA8a�g.�nk�E6�42S�4�U���%*hG|�R?Bn�l�AE �5����}�4ޏ�E�C!�)��t�>H����..|��_�L�P_�̀���}9\H<�%`�����n��i��ޟ�����$��Jl��\E�������|����ŗ��|�M��\�s[�r�:��rS�X��C��}��7����� D�cJ�{���'�
L�B]�^����6~�E�-_	�]'���� ��:������/*��{��<3c�[��b^|qP����π�m!�;�12�gm�ʕ#Nh��ҩڙ�e�ǜɷH�f�$i�@��NEU�M�%��<�R~^[.��X�y�`͌���w��;�}jkúm��m@��"�3͛u۫�:B��E<�`�y ؒ��R 'u�Y�j�hX��0eJ5��oI��fzs�@���	}����5��R���C[�X�I;��1N��u��������K�8�h��:��Wq}%�<�7m���)#�nl"���{�"dH�D;�HzU���A��L�}���Z��KYN�z����/�AA {&c��@)9�f�S�:�ŭ�	���B�}������(H����&�7yB<̬��T�-��t=���~>�p��&K�_�˿|';������M	6E;�{�F��ߥ��2��`S+�5?Es������R�*ėp"Q�p�+��(�a�3���X���J� ��2�q5a&Y���3�ĵXt5f���E|6^�oF�x�'���q��L��[���v��/O�vq��e�%;й�ϫ�<A�s�	 ��լ�v#,]q�����ka��a �Â��g ����c^���n?�K`��(�R��x0~Td8-��I���a
TFӮg��:�+��ۏ�f9��Nt����	�ʞ�����V�c�+��50�={Ȃ$�2&;'!߳E��r
���J)2܄`�iQ;��J|{11����`` g-��i���
g��x��&8�_h�@n�R'����|'7O&q�8I��ʫ�)�ӷ��G�vAWȣ��%b�!��_���%���@BO$B*����d$�*w�i%&@��EGw��W�KR�t���LTW���M��mT��:� �D󥥐l�8Sek�q�V���p��B+s�������]j9���S����B� `��j�&�5�x�������0j�Ai->��ܩ�S�f6l���l݇��Q J|g�������.�}J�z�"��ơZ;�ъ�`��_���s�=��PQ�n�4Z�e�+9�ٚP�ŀ���t�h��:9E(*j��҆/�\�{�$|T=�w���%$���w\��m�\Z�
�><7��*�ᾆgi��zѕ.y�m���Q�S~����������W�{M�K���z���kB�ꛘtgM�mƌ����K�`���>t�6�*V����lq�P�D5�ft���M�����xG�rA����AN�m_Q�������}!$���,r��L	�3F�'M�D���(�%f�"�Y�h���)�����U�6vT�-C=�.��t1�KA���O ꗖ.t��O�`��	�ψ�ު�>@u���٠8N270���|3c��|��W_��/�ep���]�pᰑ�LHU;�]�Q`fT[���HN���h��*��bP��Fg��'=h�S�-��O�4�L;�N��}���yF^`i�/�5T�wb=�ܑ8�ʦ�!���  ��~�v7|*g������=ڳ黖�u_�V����Y�8[�=Z<�k��X3\�
}Eu4��o�U��2�I�K�db��$X�U�t��8����u�"o��}x�~����Bì����p� W�D�Ҝf��������PGL�ɒbG�_g���72��%��,v�YҖ�5�ܲn�,������b�/c��0f��I�aX�����H��Π�-�&O>y�����-�.-m�7?��8hl�N����7c%�Ԫxa����!��m }����	��F���2�ެj^�����TI�!-|q+�;�?圔�Ռ`�c����J��4v�������I�~�BN��'T��6��T'�C����LK{����~����|�+�scQ�t�XF��gϐ�H˅��a�$��l;����GUPZc�H����9�GH�!�T���EvNǤx_Z�gC�l��.<�g���D���㬀�ƀ뿜s�� �n�_�f�W~o�,Xb6�쿬���X���+�v��	s|� ��_H��Dg����%*�]/��<L渑���aR��X���U꼶����=��c��@�}g�(u|�2p���n��|+j��q����3�!&��Sw�Z�0�Ӷ�rHH0j����G��h�fm��TK��>r��8�A���g�rm��ތr�
��M)���*/��5�^61�}K�GG}H�b��~g^�<�%��db��
�:��#�;#MSn��9���K��UӤ﨩�d�M ��X�9�\rk����h�f�ؕ�IU�d���#�ĊB�'�����:���Z�����n܇ʃ߯+�N��IF���PGq��Z�b*�(roKc������|���q�6p�2���;q=��┼snGK�>�{q����?�/Ho��Q[\[V���nyj|#�hDcj����C�
헁��W[Q�kB<��6K9�i���O�n�D��F��aX$��:}|�؆dG"y4;��`��Z{)�J�+V�eka3�w��h0�)1�X�֔����[{�v�Lfz��~��Kw�q��~֔{.��c�1�����=�y�yC=��qA��&W���e4��{,7rYQH}���,��T'���,�_��IV�1�%@���˭+���^�Hɰ�n�-c,��#ǩ:ʟs'TEp����)�\�*�ёU�,�<�lY|���Qb���\����I��J�X~v��$���x)Od>`���0 ���ȸb;�jFAJN_}��Z. ��J��ڻ+�H���'t��&?Y�z���Q�X�3�ۊ!�!i�O>���P���W�c���N�'��Z���0s�ư�^H �LB
��Rx�|�,�I@�A��-mg(I��G�ޱ�۲E:�$+A�!+��u|�N�Mm]�F���I�~�$+�Oh �{�@OS�:bK\@���v-��$T��g�9�W���|����^a��,�����D�^�G���,�/u�}����H�O6��������A�9]�� ��b�R�(�w*��e�����D�V��|���ZqV\�z����hs�<��V�>*SP�h��K뎶���Q6��?�}0g�����N��C(U�*�H֝�5�?���f�*3��8Y��,�jCX�ؙ�#hņ���{K�2�����Ww�*z�o1�ּ�]3q���g71�L�a�'$�^��x�\�����-zP{��㶷��js�Id7J�p�#�c�<����:$EI��:Ю~�� F�=����lE� g$f�%YC��<vy
�>���Y;�>�Z=����$������VZ����a��Pޯ8�����^h:(��R�����4��ؾ$���<2#("D*�!Ҩ3���XĖ��0�촽8u�k0f"(�/v��{�l�)F�>uС��+���'|���!��V�W�Q�
+"���,�DnJ.ԙ� ��0��3b~���.'�[|�o��;c���ZM�6���ꤲc��h�c�}+�
�����e�*8шI$k���]�Z��1�������i}��N������ުw�h��
�Sd+��r����1
�~ �޷H��.HX��pd�mY�ч���)�'��*�0�j�d�����r���i�M݂��aٴil��F����
2��J�Ĉ�
�����
�J@Gw��x��T�X�{�����`;��7 ������{�V�H��x�уd��J� �Kk�"�
ÿ��7ƙδ�����0u�Xnb�g�2"��h���M#��P���o�V����ޚE[B���_����-�u|�m�
a["�������V���s��(:� �E�}r�2���ʜ��j�5��@� s#os��f�F�`�k~�\��/�����N�L\}K~�HA���˰m1�`U+�q���^��w�{>sY�i3���vK���0��וWHS���LkV��oFB���7�=x�d�����	�U�9# �q��JĈ��_�(��
o	;�����z�Z�3����]F�h��%`�ZoF��{��tg��jX�z�!s�z\�C�f0kr7{��,�g2I�]K�qm����C�w��W��#������П��"�[ֵ�1>�v�N�nS�����
-{%��W7�����c������}G�V�v�(S�I�ٛ�������P��}��~V�(��sٳ���'��i'	�e��g`l�#c#p� CYYd�"�|��s�����K ;~]F���fґO5�/���㾬��L��R!VY^a,�em}�?wC|�e �{q�k�{P�Ză�"R�[������8]_����H��L�q2$Tu6af�ok��ii?`�"�n���\ݤ ..a���Y_ߓ2W02�[��Lk r�Tz�J��Y��4vl0���.X�����\�Z�ri���U��3Ȋ�UBg��|�T��8��0���}*��}�������N-�w~�	�M��wFc6�����{��J���:��~:��������bOȠR��f�:.L/p�F�tI�˳�Y�~������m�W�"�6Ctn� /�Z��J�A��g���S�y� ���>_�}�UУpӣ���p i�Ѽ
Q��l0�7c��BǬ�!�x�Fy��eus�c��՚R��k�dt�$��6R�+4Ujǣ��b=���c ҸM�,��AJ��˂-�(��^S���Rn�q3����%�1�W�w�2G�V�,�w�"m.�~�{�)Z$�S�Nw9��>�,vz��*��	�g_���1o*��WFF�x__̇����Vq���=�4G2�R���w��a�4"��'g
�L�������Ԑ��bA���	x�0h��n@5H�������	�[����|�2��_j�f��ayY�3��T�7�B�D.(�Y��[QҢ�ތcА�{YS�o�d*a0��l����^�F�>X��9�Hr)�+l�$D�d��n����d�
!ӻ����.RG�\i��#�1l�(���^fq@���>��������3�m����3�-�+���
x"j�"�|���6a����pc<ɳV(E����~��C�Ĕ������ �8!S�!�z7�ЄS|��y��K�ۢ���Bw7d�e��&^�f������c>*�Cg��##=O�D�3Qq�qf��Ɔ�Ơ=�cQ�_�iHR~�������ܫ���������x����N�4�\��9�Q�pj(�c��d'痒+;IrT,�눣��1Y3�_?Ր��~�"�L��F�IK����Rn���hGyn����dW���b�N����&���̜`R�͕�=b��U��*��v��ʦ�!�׺��}xU�ݍ�����h�7'{p+NKw��9�`ث���Uc��2`�g�I^ݱ1�A��<?�U�%�;NP��0���M ���e�����&����lTNG��Z��m�t�	�� �+�ᬜ��9v�5WH��>sR���rNլ�&ok��@<� 8��lsd��t�aX����*v�>��Sa7� k^:�aR�1�IUs��7J�St���L	� ���T��J���˞U���[� ���Q�v������,�8^�6�)�2]A��A���
E�	�?@�orY��4|wÝ/2��-s���������Q�gN�иX.�$�y(l9�׭T>�Q��S���0��3��pZ}y;XU�%��Nt8}y:��&��}��]��0����Ԕ�&M�9<I-J�-ץ�j8,u1�u�L^�����m�����[5dX5	�S�?#�[L�@�&�T"4=��?��5�V�nVF��K��=;�j�#]	>r�D͙bQ�r�i������kt��_�su��H#1{J*�߀ I�����JE��$���[��C���ٔ�4�p8�rS�ZQ����Z=�m���؋�l'� t�=�谒���N
d��R�6���1<^
�K&���`y
���3��Ͻ�(�&h���o�1�(28��˿�ƈ�u�@�n�*9/����v85���Q�io,x��)fj����D�=�~3Q ña��A���A�_A].H�6��nw��O�~�h8��F)m��Q��>2��܉u]ӳ������"�j�Y���4�)�[)n�W��>�vXb��k�j{�e�H6���H�{Id��Q�;[[��ejW��:��0tʹ��=̍[�a:�`�7\�|/��O5ѭ81��QP(ǰoU�+���a�_
�@�vE0��+�s�K�8|	PP�'��,͖xq��~P���Vz�[ ~|U|�7ڛ&�Zh�#�M��
��9\�D�ð��s�6>�-X���(�08�I�v�I�!�oAU}Ӑ=���_3������:iګM��c�ė�ޣ�峭�[��5c�S_DWy��LM9��_8�AmKH	xHka ;�D��h��ZT�� i��5_o�XR�R�e��&���1�[��o��6������\|x�"{��I*@��Zr��!�h��a*@�!���� �^r��P#zCm�[-��㺐౹4:/
λf��j��|6�t:�R�!�ٕW ?��Q�a�倪i�Y���y��D$����ٰ��?bwJrƥ�ve�LI�Qq2E�`�����"V�n�Fi��Ze<{\� ڙ�[�}���X��!��ǎ�:Q�eՈQ��&g�:	"�²|)@���i�X0�іц�b��'�:�re�����}�p�?��s  XУ	PG�<Հ�Y�7qŏ��v;�a�m,�j_̚{}CFSi-MR����������˒ n��oǤ���Wy�2�w���u��̜>�{r-�B�%mn	 ��\�� g���|(�	���yM]Q]��\��M�7�y��S��$XDĊ{�$ӗ{�Bչ9�!����T�� ���B�T�5�����'�O����ǖx�ks���{(/C\\�;�(�`�x]$���x\(��g��lg~�M���'����c���ඏ%S�Po?��1uk���k���.���@K����_ܤ������B
w�4x
#x�������������h������0D�Y���U��\i���q����9EdU����9xk)��j��9Z�lYw��U�d�GL��.#t�t��u_<Ǘ�b�A�rsLyv+���Ѫ�pSZ0ki����M�I0��R#��D�H��C	���kۍ)XT��.��Q���O}߱���5ScF�u)MٮAM�w���O9�פ�cų��<-�l�����r�Y�{x���o�� ���]�x���Ld$�`=�G����*<];��p�&C�2�6 �����J�j���ἔ������8��2��˅e� �"0���$��J��ߐf�H�}p�y�M�r���pV�9��RR"�R���Dj�T�I�	��ڻ��3n�M�s�Q�;�2�f�2;(��;��w�z�"����JK:'������߈���}O�1�=�𤩟g�Vb5�s<�=ľҧUb����|M���2p��R�g��T���j�^;�k�i�sxQ��Pyn�E"��5��&5�%U��fm����Hg`�}�0��2�~��M�(<^͙���-��FGd��&ք�Z�9."ګB�
~���?��Jn/#���jK����ח�}�`K�-$�a��J�{]�p�E��w�v�zZ�j�+&���F� |���f�T>��򮾅<�� ��_4P�Y��7������,�y������q5��z���˒U\�թ��VK���񳅼`
�*��?־�ɦ�PL���At҂4�r�mVe>gh�Za����iɟ����@*LOPy-�$5��M����F���ك)W"��b�O,{�ӂ]*��*��<󒩊eN��3�@����nE��Fd�͋��Sʍ����F!,���0%��;��".�q͔i����&[8m]��
x�Dg�z���% ]2����$���P���B�#t� ���ا]���u�����U#��c}{��=ǰ��sb�V]�r��|v5�/�����v�z�����dD�*��� ���T`��d��&��}�{'Q���u� f�5�5�Zq�߉nR�]d�p�h�.������\Tܾ�Y`�e�/�GT �ͬw(o �ea��p��{Zߖٴ����m��� ���ͤǈ�Q��0n�n�Tf�B��8Mh{���vG^����識VB�h�}������t�y���#���2�#�rG�!J�F�~%1���f�g(	�k�~��
�zǳh�����
�8j!�t���d������]7u���&������VT�B�e�=��SV^҆�<?d�U�d��X����g�y��fΎFw�jo7�-�z�s�\�?X�ɀ��s��.6c9��f$J!�Z8�H~�p�Mڐ�L!��� S5s�*�2�O
+�=�R>�N��3���}����=�-�3�mm�SS��}�gz{��u��:;��_y�z�wDb=���=�fYS���A�Ň�S�/�/���Z����dl	ށ<yY���*��\o'�r��D�J1"j��he���_jh��n��䄷t���B�N���P���aT��r�P��
���݆s����ԍ�]�q(������a`�E��)|�� ֆ�T�6M�^�� `�O+(s���ph��аD&���6�m��`��fOZ��[���wa��ȑ�u�����8�^����������W�X�8��'��������ϻ,����8�Z���O  Fɯ����c���5}BH�@mY�'��u>sk�B(��7�.��T�|ݻJ�����}�A��4��A��i��).����eo$/����F�*�5�_X�R؞����\�������{���f-�����.W�[�*<[�){�J��Ll�}�⧎���Yk�7��r�����8\�_iI�r`�Ac)w�$MR�u�LI��꧋�1���_�m����'��0�`^CĔ%���%w�Sz0�k��,-�6��,��}��ҋ��lBn�o����z+R�%S�DfX.��	D��P��W�r�4k�4�#�У��zT^���`���(���0z1�Z������	J��2��Y,�k�I&rG���N�����=<v)�ffj����W.#��V�m����/�١fZ�
ږ����1]����{x<��%�W����Q�U�.+u7�2���9�����9�-�� ��8�u\��
(����ϘP{�AO�?դ���O�.r���,��a���K���Mh��G������.i����	��M���H�l�D$���°�dH	���g���^�x��$��lr�����-0󬾒-�U	�R?[�{���ܮj~(��dt�}�@:Wz�g�w|@��@��<rr��?����vY�,� u������n�va0\�����%�������+�f�mZ����	+Xq�'GQ�`�m󡗲$����5Y��cDQ����]j"'��4i*�*�_�!��������I���>V�l�R[�m���U/�տ��J����I}�`Z�ɽ�_�i ����R�쓂�K� =|���D(�;��'�M/�sQ����Vj����X�L��ֻ�] B�42=�^��>	�U_����p��5/�-K��a��9)b)��	vo%D�����]�Z�æ�ƅ�N[�O[�����=�Z�����K ����k�qG�y�vٌ���0�t�[���r���`�M(�#��>KX��Q�C+VB-E��E"��U#8��?!Mpv�~���8��	Q��0����hVģ��)T:RSd?�z#�VwA����ÝG��X8���&�{���I�`ӹ[��/x�%��l&ܖ�?vl��qR���D��`g�sc����Q�����gt�b+��e���ԩ�!� X�Ƌ qZG�2�4@u�Һp�����Z�i������	���"��qw#�t�Z��hi@B4{�_����R�A�O�4���E��	��(4��?a^r��B���\�,l�}H��9�f���7���~�Ys_��Q:k�U�ُ}}��TH�F@�P&���;~?TN���-��s^����Ejܴ��I��}�њ�������K`��|�,��sl��0��P�ڏ�Mw��m�=O�5��Y�X��dy A��=�aܚWZ�#��4���K��s�v��$��[�e���%�E�+��R�SN�1�6��Ґ�5ۉ�i-rz}�٢h�"t@�ٝ)g�/���ڦg��$/�7����Y}r0�_��7�&Dm�<�.�S=U�@�5x�ݍ����b�aPL�E�͑]�5����R���X�|�³4���&h�q��.w�N��b����g�P-�c��(L����}��c����T��ɦb�� �G�}�n%�3ZP�����}{�~�(�ԋ計F���}�~��K?���_�ʫ���L�ܗ@�?_O�����򽹭��=J�_�8�QK�/ �"�Z�� )�0~�L��؅�O�*b�&�x��lm�C���XX�rg6?�nZ����4֙Aab8?�`EN�<�H�����7��J��o����9�ˤ��'00��sU8�N�L�ǃ{xӋ^lR'��y�ɼ�k�QY0;���y�����չ�!��4k�u�i<.�J���8�m鬋�	$��^�@����ky[.�-�W�>Yz��F>����~ �%�k�1��[˿i ���`����U��1gИbi�@�2����6�\������肋�������)��ˍ��A�7Lh3�3�}���?�s��zϼ���ȱ1����`|�����RK�(;"��*�D>n�ki����Z��pd�{�і-��׶�W(��H��N��(d�6��+�uq"8� c"��l������z&�#��E}�$A�3��l*�UabӰ�U���4���>R_w�^z{��ɥ��햁}�er���&����6:��7���Mx���C��0�4�(�i��	Bχ�Q��z1�6˃ux��ÌU�=�כ��k �6�Jk\ϐ�d���Agge,�*���_H��������=��I'���^Y��ݚ�#�C��ѡZ�@ͧc������O���n��z$e��=����/�\d"I����Hnܛ[nA�����ף�7}	�俈�lU�j��.)��y]V�|Rs��97P|�6��9��\c�����0�B���C�D��"��VDk��YJ����l�"�^u�86�l@�ĻS�>_�����?M��x[�|q���&��Xh�	�QLo��ą"��aϾ�0�o���r�*� ��<IU�1��"�#�:�-ۖ��d��D�t/��OuE���>y`���Z�������^�(rӊ�~ƿ`v�F��]�����M�V����V>\]�Wm@H$x�0z�'ꂾ�r��ўa�P�S�*�Ct��q}���]>����LB��	�¨�hhrKL�@�����WS���g�C�#w{�WT�S�=S���%\M����7�dNp��x��)���5Jq&O`�_�I���B(���-�݃ǀ�yQ4�n8o����u#,ӟ�½��-T��V#.?��Uyz�\�=y�˹W��̟r=��N�;�ɺ�8�P���@ox�:l�6J�^~{olC���,�I�<b$�){BI��Wϗn��@��1p�i��ں�&��f��&}�!��w<�Դ�S�FŻ�)��-⤃�d��$��`A��w�p��Lç̓n�,�#�b��trb�ܜJ��빶� ��E��rK�� KOQ����F$�Q7�U/�,���&�M�@���I9r�Z�{`����T@�EE��ԥ��iP���ah߳S�Q���H�1�?���P��2R;ȱ�[l�0���wO�փe�������V���`���E�^Sǖ�������{�җ��Z6�$$���a(fGN��ێMd7f�?���oE�9{롌�~$���c�f�_�����}���X�K{
9h�2dd�c�2LDӵ?<�����1�~���օ��4��
���w��T�����u�ٮ��ɒ��w��	<���2EǸO��~��Q�MAN���x�=��zO�&Q�d��6��dl���,��*�Gg��t�9�H50A�����{m}Hh�;|�D)��x��l$<Q+�G��}e�T�4�u������Ҭ�o�G	�iz�:�y0�Ʌ�u�ސ��ϫ�O�m�<�Q�?oA�3�%���t&D�cڻ��,3&"!����?��E����;�֘"%|7��`�ۻ���6o�hG9����:���g4&���d������_��N��#�&5d�����7&O�� ��M�}��0���'�/�v��,���S�a#:81�H���#�Q�����6`v6��~K�)ף�������UE1y���Œ.�@�G�$W��BSg�gU3p�����(y��_�9 ?�}nV�7����\*jz7V,H��\�Ď��+�iDdq)�Iy�����Nv*\�Cs���tp���@����_r�,7��{|�@����/�zqMh�L ��8�u���^�<b����w��� �+�>FS�!+�>��f!��~$�cIȌ}߫�n&j��6������o������o8�	�rP07�	���m	�z2L@����R��i���Dvrt?OӀ�ɣb�时q�s��ɔ��u"�l���Cӎ���6���R��@Zz�ƀ�q��GƏ�P�Q�Pfwε>���{��Fj���p����s96�82�y�\:��C�֚����}���>�4��r��qd�d���/�5��	I$T-�m�;���+������4PIg"���<2�P��m��ٹW�,\���砸��_�����i����INa+��Ȯ��h5��X��3���]�b�Z��^b�wL�d�"W+շ�^���������}5=����h�݇t�,Z��D�pi�(��*��f�5��)Ŋ���@8�{ ��r�6���Er�.A�
����<v�c�*B�8��"o��{FW�m?v��Bo`�J�B�Z�Wh��?���g	 k��@��ۍZ���I�!�T��Cԋ�'P{��ߖy����� ���w����8�ii���=%�78���Hs��^����=�'�/w�-�N0$��{�Ȋu��E����]�,�qWn)2�%�qJ$k{�����i9Ҭ�iրi��m��V��Gh���*,�=I:F5ڜ��EҞ��DFy��o^��)����^��O����jp��R8��4�P���ViF�P��|�~��q'�遲9�7dn� }D��R8�>���ۻӄ��'��O�v݃�-�D�!\芚�@��K�J�-|�P��-�<|;p.D�g+]�B�-�Z�cp�	C�=���1�<cNB����^J�i�g���uk0��6h���	�#��LĬ.�ٰn�E����
�x0]{b$-S���k�Q�<R�
���7��!m�1:,�:1�b� ���b�������ƽ{�d=������):3�Jr�(���t�����\�D �
h���ya�c��d��������w��g@����d}1�W9���i�p=s�;-l����,���J��`��#>��zo��n���e�RJچDTt���s�F�8~��>�,{W�F������"��'fp}a!|�-�o��ީ�~(O�/iK�э��2d5��^��67�����!7N�勁��	)��#4���4��W�V���5!����w ��$����H0�G_Z`L:l��?�Z�^,(.�!�ȸ�'��z+^Qi��0�*�v�2�q�w=[��4u�1�"�͈�ݱy%j�N ��43"Z<����k�"��"�g����ǏMO����%�0˂>So ����[P�n�����L�H�� j���@�U���G+v��V0��nx���J��<���dV�%1�����Q>+�)(���.�S|�G2Å��)���Ѩ�J���ჲ���?\D� o�4��*B��H�. ��ͯ>�L�I��d�Y�O=�'SB]A�ۯĵ�QO�ob3���?+%������r{�����8E(d�~,ۧ�	1g�N�V�����Q
�E6�S:	���v�F���1ا&�����$<hQRV��Nm�|4�d��:�2q��X�!W��~��,�p�����a|��*6]�C0��,S�1���GY�p��8<������^O�������]��f���A^E��Q�(o��AʟG�c��>"�<#^f�~!h��gY<N5����R]�S%�н8R�U՚!fF[s*lY���l
;/��ލ��&�@�����tGL����E�L'�UZ���>�}��[x����)y7�Z`�*�
F�U�`$�Ǜ��yf����
U�}�-�R�?>h��<�c*|������Ѡb��g�S�«u�GԻ)[]�e��L�e�X�䎮�W�+������9m3���`3��h�Vʯ=,0����x��nV�=��Jb ���ֽc�S(c4�Ue�%��%]��c���L�r��B�$h��1am�4�G��}�ב9O��P.� wa�X!_$s���	���v꾆=��b�/����,:W�'��6�Y���)�V����3GU]4�knT�)
�l��u��{}��ʰ�ϛ�ɍ��JM���h8��-�D�������8!��h��x!������[�>�Z������ÔbN��{�fh<�3���9:��H9W_�D��?I�9#,�U�h8�HsV`&�=G����`�>�t����8����Ed���4��
o�R�L	�+��#1_SN�Rt�l.z��ϛ�j���EhZ|)8"D�^�4��[���ɇ�^��l�c���w�4R�y��B�����YO  
�5ƺ"W��8���@FhƯ�ҟT�����Ȱ����γpW����8+�(LǶ�N�e	Dk�~ک�����aa�T��2���,z�'����˘���?ը-��MN{v�J-}v5q�O�n|̌ӫoj1F3C�Iߓ���������x�k�S/�^�, N~���y�Y�~�@�u8����/��"��!�����)�Lg G*��3�p1�Dт����Y4�� W^���s�Q8�"a�d�T��q�Q�B�tlH���kأ��s!�n��֟>L�� Hz���鑹fm��)ezme��al�j	�WG�ɖl2�����V�8�̗IsrJ���>\�z��z�}�C��r�`�)�/��Ht�+����(D̆�8���4�)�����:���xs���d����Ƭm�A����;i٬ą��K�f�R� �
ѵp��ǰ�����OE�y���������W_ߎ�(i�N�3���/�z꼧�6C.� �)>��N���kc��;�(�x��?�x]@|u�9Ѧ��v:K ����g���wh�k�SZ�3:�'뾾ٜ<I�9�ku1�Q4H͡
�h��re���<��U�o��ꀢa◁\;E�)����^��Aزa�W��P4C�rv�ۜQ?�.��	BZ��A�����zRT�hi�.SE0�![���\-�-��%�P"A�Y������!x��wU{�Hɞ�3Zh�d���.�Yf��vA�;�*��Od��_i�z��0��(�y���Ӱ�XU���ݯY��Qk��x�s��D�G�I�����F�9+�OT�sv�6�� e{g���y�\v��"�B���Dw��7��d���ڂ)�	A�:�h�������i�j�&���r(ck�Ď�R�_F�c�:��S�{��Lm�YJ�y�{/,�ש�'�+�=#�r�_J��1����F�5<�t�	uA����@
&��Si�nF�����=4��x)kZ��ִ�ˑȶ�$K�f��]�0�8)���XE�~).�&���Z��X�4��:�^1���'E��p}J֯� D��Ar%ݢ�Q��:ѴA��n�A��,������Ӧ�1h'�x�	�lc�&�TEZl�r�
kBe�,����1K����yp"T��<x��B��|E�\D8G��@�?���Z�\p>g���t�Uv���l*d>.�R	 qTT�|~V����p�-��j�<\�1B�k8��&��2˵`������CL3�_( B���;�'�N���l/e��u�WJҹU�vFj4��Q&6�X6�GgT��´��Vu�ƚ�2$լ�a���� ��WZ��o���.B��^�'������wMg�9�͢f��):�^���I��F_��,[����L�3��m���l��&?)Kս0A�X�˜Ća�>u�.`��l3��y���w�a]�F������6�K�������06m�>Uǘ>*.z~� �PV�$v�Y������`S��	�N�?�Q��{�N�tI��h�W�G�yD�Xv�l�g��#�ߓ��#��W�M}�gK:h3��5W��S�M�R@z)lj��4R�U��/zuz�*�Q����|����EE�P-�8f�F;�0e�CP�ީ�ia)���9�r(����IW����g'�y�J�(�A5i�
ۣ�7�ˀSGi�eH^|�Ӕ�����U h�����)i�2Ԍ޿=2�`A�k���s:���{s9f� �`��F�=e6z�H���%��ʟ�U�$��;X�@�a���`%��st�I�w�KI�mOj���N�0�0�R��_�%���(�c�����Mf�Ϊ� �ކ��{�ec���K"�0�Q�OU���:6[�:� u<`�R�S���}������ı�>��ۄo�����E�\I�7��ض��u���T6�O�lHb��y���I?C|�GA��XPY����E��G��.�z���TA����L5j��<�Z(�'��g�>1\��8zP/�6�E����$v�D]��)q�����_D���o�%�U�'�
��v:G�Xa�G�F�m�3D�M�{���}z��G9"����C�Р���K��y��T�ޫ���Dnڟ�7T+���.0[Vw�N_��7]q�y�����Q�_Z��AY�/�9l)d���@�&��2�r��r��$^x��+z�m�XO&�-�R�w��U����$�H�	\_�}3��鰘��c�j�����9�l�*ǟ K���Bl��V}X(����S4�߽Wj��EN�#��2��8��.4���M��"�s�-Y���	�4k�|�>�K�����_XD\�wj�x�9pUE��%���>��@͈�z &{vy'<�d���uʳ�.�3~e	�t�Sd������
�2C:#m��.�����;����q�R�r~ZGr@�<o��n�<�N�{��册&b�TK]ElBE����������[<���٫x7�ՖG�*i���W����-��D����4y��Q�[��B��^���q���Q+>�R���k�&/�G�y�@f��M	BoF��0��qCGs�3���6�]3{�����ބ�8��澞aĠ-��|�eaH��[�-|b:��1�c4�l)9�G@o#{����4-�U▧�_ӛV{:�C�������aE�n���C[����zkh��Ѥz��E��ms܃���]�(�q��7����]
�J�_fTl9Sq`���
��hsW�?��O	r̋g��9��<?D���zVD��ջ�?S��eȒ�4�R��x��x�̤�D���hh�̼���W�*v��4�����y���DE�hL�D�������H	U��RP�� �$�D�N���P�#fق�jA*��3F��J#_f�� �M|2z��Q��K/!@:E_<�3�#z_T)#׈�Eݻ!Ə����khd7H:�u^k<B�&Qy"-_F��(����&�ۅW�$
˲���Å,*��@⛨�R�(��pz���"�	,�_�i���}>�p7�㓝��*�G�A�;+�2k���!,.<�S}x�:nY���"��)�Ҥ��܎��NظO����Q%�1�8�
z�J��1zE�]rI�
�9:�&}\��L�߾,���:���^4�H�WH���\�m�kM��ϵ���O�^��M�X��TcUa�ة>;����:������X�h=�n�	b�Fó��پ�\V�N'�ȏ\1<\��92@[�h/�@0�(_ w��BP��u���4�5��3�'Xٛ[AQ;}�&���̫�i6��%B̷���k^0�F���������0��`��+��C���@g/-w��E>i�C��䎵�5�-��>W��tO��K.�C5��FP��d��Oɼ��U�O�򘄤!��)��->��Ա���.�/ęi�t=�B���B+D�^���Ԩm�Fg��5>c�}ǸE1[@��+�ː7Р��;� ��^^��$��=�7��\c<q�>-�C4aZ��:\����>�J���x���䝾�a��i��j*��5No��2�s�O�T������Jw��2/��UQ&�m��\M�� �#ô@�i�NqV�	<?�7jֻ�H Qe>0�:��9e�Hkx����
{��/�S��7`��=�� �nA_cc���'�Pݞ�9��Op�}�K�b=PG"T��t���)�5s�X)�(>R��c6�B2!J�֝t+���=lǪ��O�������p̝��Zkft捺:A�x�2������d�1�7����O_�4��y����HK+��)�j�+;��\8�2�#�o�j��]y�Ӳkxx�|�,Z*�e���e����dwFNˬ������R�w����r�\s�\���P�]>o���F�`xR���=_��o ��L��2�`�'�t*��cf�{v�)T@�ɛ�juRN��_��f���r�8�H���Nq���FO?��'�{�nFM�I�Cļ>��P� �KQ�@#�$'+��N[��C���90��Ňuh�W2Tr������������qG�c�� ��b�pÄ-_����� ��/+� �2���g�����k	�Ρmu$ݿ{�C<ԢB��cK�_��Z�&3�Ƒfa����ZD�|�Զ�$ ��V�O����="�d�n�H
p�A���0l��h�o_ƚ�S,_k�D�h����6+���;2�fC�@ML�|D�m*��s�z�%�g��g�ӎQ��8��e��gG�%G�ފ��1�W+���y��^rSiD���׽
�L-0l�ATa���zU����4l�f�J(8~�مz6��E�5Qz�7[��Ṫ+�iC��q��I��!;�G�Z/jĿ^��v[RVr���a�p�Th�#<�H#�J�B?o��d2�4y@-�5�V������+%7�e�	[��vԆ���{Q�x�#�\p�i�h|\��~����,��[���'KE?��p���14���?����S�W1 a��5h�Z�W�X��QM�Fͯ;*�����>A��{�⍪s�����t^F��U��%��N�[/hCF�pc*��Ni<���3�~�ZY�88>[�Ҷw�I�S�����jX��+�+��g2��^��d� �(P�~4O0�)����V?�2��̰RQ���ɇi���G����%�Y�c��C���'��g�G+)��^�|�̃�(�+iM�|2��_����xf��)�X�D�Y�P���m�Z�
0�x����B�-`Y�&A-�w?R$M`P���>d$��\�0�Q���9�v�!,�+{��GG(�G2?R�t���[�c�fE�Ĝ��kV�ox�b��U�'�Q�U�gᘚ��h�l��������g������"1.���u��Dm�7@i�EכƑF���m��=��ѻ�U���O�$��V���I�PTu�%φY'd1=�M�;�Z��#7d�6!��`���W�����q�%tB��g�bz�G�g�`@��k��]0Đ�QI*jA�G�\�kX>���o��´�հЖY��+��N:i��,��  N�[�X�U9'�͋f����4���f.bQa�����Uws�a�<!"[z��`��C��m.�K��x�QxikZ��řm����y��g>|st�7��]k8Q�T�,�����	��2�ٔ^I�l �F�.����	Wd�����nN��l�lGf��u[����b�󙳊��j�/���'�TA &��&�������%I�b35rӐ۾����뚅INC�u0�{U���R+̖PT,�XSL�Kxٛ�1���	`��"s�`�r���6�b�!�$�6+�HNH��> Vhu�r0S���G���%)�����}�0f����V�M�\�����ma��G���;����Q�� �^"�0
O�~�=�Kp���z�]ph��@������\(�����v��M��p�q�x�%��~�Ҋ��^&��U���cx,'�<��ߴ<h��(9,*�
ZU��F�sk�II0��n&�b|ݼR�姕�7���\�I��O�;~����m�7�eI�8@�)a�J�Q�)G���A��t���K�=ǈ��Pf��6q�De���@8�߇�6�m|T,K�u�I�ėšY�	�����7Ҭ���^�I�C���4S��8�hwBp[0)?n���؅I�o�vY�]��V�����c)9�E�#�L��IN4�݆��t"����Jϡ�[�UH��N���-�\d��8ή���Ktp���_�pBB��'+�Dŗڡ:��8��EZ.e	���&|�W��y�l��R�45YM�S,���G��S����aC�`�91;����s�� \�!,�U]yJ�,�Y���}�*8.���,N�(2�xa9����h%'W\	Y7u�oXȍَO��3:{�����O
"͙ns�:޳��[�`�5��MjD�����,��T
�{y4���q���C�E�aĊ� �.9���s'H�gn@)7rN�es>;LpΈ��|�3�U�����	�LU�Y�av4UKx9�wV�WG[{��#�}���SS�68�e�� B�]o��rl$C����I�`OJ��j�� �B~��pՙ�B�u��� �\jc��nS�����pTH�5� �Mw�^�"����r�O�++>��z���&�C�����/��y{K��P�$YӇ��W֕so���mG��J��hۊ�4�q��P }旁��d< �M�h�|)qX(cx�#�}�"��5&��`��*˟`Z�<�[�;�<�5�u�-��W��1sXA�Ǘ�gb�u���F�g���;�*T����PNPNAG��p%�T�����׹��`P�������澖�}��0��K)ɡ�ļbUcT���ᰌq_�m�	��i��m$�B�1�{)5���ۺ;}��"�/ۛ�/�s��8�Pg*�gJ��e�WEB�U�(�"X�z����!������/&s=�ų���V�Qny���ߞ�-�VBz0�(��l�����G|�A�{|گ�׃:BJP�W<5��'x؀�-0^�44X�UV�vQ�#��18:�@$���F׳cq�l�1c�d�h\���V���Dt��;��!�v)-P)��m&�n����h��ЦpO�>�1)~�a����,�m�	�(�I�r@j�u�QZ�2Ɏ�������SL�eq��I�7.�haK�ly�p������10[HZu�l�
IRJ��u��k��f3����h���P�9�D��֏2��?�w�ڒ���>��}�ѡ��)�gF�����9�H1/�ȕ�9&��o��Y (��F��:f:�K_�@���9[o�/�P-ڞM_�,�2s���ن��+x�'܀<܋��c�a.Ҧ�g��+t�J#���M��{5c�:�*2kU:f}����2���j��h�Y����%���ؽ��v,��*n�m�Kf��'o��VR³(�|�z��E��ؒ�Ά�!����$�E��G��*��g��t��w��\X �Ҋ�Y��L�ڈ�6؁��M��7�f����I����T���e{�y�t�_�_���:�¨��nH�vB���TU+�U���o��o���(ur� 6Y���r���p <3�U�I���w:J�����9�6d��t6	ޔ��|:*6�H<�(��ڛo$��Q���xyg�I�����bȷ�[q"w%��	vuݔ�[뒾kDY w[�)�����M�U�D[�T��2�c�0�)꼎����Qt�j��������okpu�]�sL�vO���CW�����b(̴y��K`�-tf����ɻB5"�C���.�m,�����<(�%&�#���.��N�%*�O�ߗ���:њ�@��H��ƍ��y1D�:۱C��⬞�|�!�ˈ����nv1Sa��hCK� �եAQ/��	��G0NG�,4�Z�%JM�i��
|�h0�����݈�#���t��u���T+�o�L	C�!���H����v�����u���k�b���e��q2-oT����n9���ݪ�@O�H�}�T�U�S�������$�����{����V
��1�֗����h���cu���D��Ƅ��N�t�Rgdd�&ߧqt�[�f����/l���H���m�)p࢖{Va�cF
��q��_3���)�v�۾ ,����V<g\�w���Ċ�#�<"�2�X�7D�(��`(�3[�,f"iO�Jg�)"�r�ib��@d-Q�
$�^���V��p�=��#Y��w"�B��hb�Š�r�]���Z�����X$�
�*�j@0L�HB��V<������[��n���yQA�x�a�G8�+>�Ѓ3�8HY��:��\A���GkS k�^TY���"H��4M�ˍd����Z�����2{�5?�(藅[=@�E��1tS�4x������@%s������	p.�#�B �k}��.���]�r��2y5�D���w����|o۶o��S��sD��/vխ;��?6<RBu ��G��z=U�j�������I�ztM5�x+����jɢ%��c���wG�UF��j�{窝b2�*~�f��{������{]��>v$�Y�[��K�R%HqJTk$��almy+��ʏ(�C��E����7�Û�㕃t�R����e����p��?�]��*�տ2f����/h�]sW$/x�ڸW��/(�ɭ_�**�E֛��Q
��6��)�\�b�I��y#-��*|LKY3N�"�#*`)V��	�����A�Z 6�,H�|Qs�U�a(M������t�0(+��m��{u�vRr~~�5*k��rHr��jO�B��u�/A�o0��p
����<�\^�������p-I:c����.n#��.5�f ����E]�N ��3�B-�\A���}��(3��fAj[�G�	�#�嫫�o�@�7�IѪ͖A��G'�=h1Q�yc�t�8`�n�K��X�|+u��Jwː�:}���48����(����M���g2F�4�%�o�oY�nT �������{-��e�+�k���U� s��B1�A���iX�t�
�U�����9A20����w7usS�#'Y��m��"�L۪�$�g`W.�D�A�Yc���:�_X�xrUշ��rX�='W�Ԓ&9IH�[��2*��բ�B��؏�ދ`���-���ͪ[Ɣ����� ��Mg���#�h��
�L�+%<�kW�t=�4g��	�s�
p�&���t�Z�`�,T�F���h=�$7@)3�6�������Y�����ZB�sL��r�`�#`�R`r�[�?n�	>q5���s�]J^�"�~�gS�3��Kh0�C�D���Yn�v��)����?�����l��Ve��C�`Z#�%�h:яo�W�0R�r�E���|L����{u��E��4w� ��^�N�A@��tX�n�!]�xCJ��f+\��
�i>�n��D6Xq~Ӱ�����+P�ۦ��x�7��E<��h	�3[T��9�/L,������X�����.xJIS�]);(!z� *n��5����R�S���-l1{1-��3����O�t���.�0	[�V��l���uo�Ϯ��;�\
�w�F9Z���l3a�2��A���>[?��g=�L���"+�?[�/㫍��/F6��?���SR��"aط��}|A�f��8. pzC����������ȡ�J����	I�b#3nZ�(�2\9�Q�s�5'~�|�j�w���B�Y+��\��vn�Kl� u��N�i�󌈰��ޒ
=�Ξ�9�)�̷G����{rNCm�]wEK4�kkЁWF���@���`e��5�	K��ȸa_稺��J�\�b����;xR�i6r,S��s��
xʶ����X��.�J�,N!�B�S��D��w��/�-" -K��:����>nb�&=|�Eau��>
تd��,|j�{�����[��ũ���($S��d��N�HX���Ps��1�'�śZv��l7O����Ǜ�����Z�zwB�$�d$V>��@�4��4��PC���KMh�|�� ��e�8�M��L�FKy���Uъ@��=WңX*���ɂ��뇺MvD/jUyLb�Ƴ����D���23>�'x���d_�����Kt�,Z/��D��܇��C�م��]�M���q�SJ|��W��6���
�Ε��}w}Kyn�E�Mk!*Lɷ%����y��73�n��\;j ��svap�֫5Q�dv�����U�#he�"��F�̰Y�$ �`�2�,�������HY��`+B�1���c��b%�k��/j�n�7/z�Pյ��/�q@��9���!{���EJk�5����s�5F���N��o��]���75YMm���+$�6�/	�����z��b��-\S��+��~
4W��1��
�A��s����0��-���)�z�"�0r�u��r�;�;u\����*�qS��}ά�;����\|���lq�b$��V�>�K�C�]����hx_��1e�E�Ym���zb��~|E���~����߹-=�4ٮۭ�>�Xߘ{�_$�����*K)�
�3v���KҺȐy;�:)�̾\CZEږ�S���
7ݛh�4>쳥r�q���ǽ-�Ōf�#�L270Ty�.��NYc��|a��b,�ȑg񙙫M��u͖-�/&��`��. ���dd����A�o�u��1�����5�����<&.�
�|�)�����gx8���V��:��6�a~��%��a�����{� i�1C��ꑍE<�8�<���ߙ������^N��7v��W�.�� 6�z"~_Fk�8ݿ��U�m�ee�#�Cz@���X�9�$��i����C%������KLZ�1B07�-d���.���"*Bn䱾�7p�m(]%�N��hCE�GM��Tj�Oո��ũ�`6u|�H+"�' �e���R��@ *whwx[�ī���`'�iNڕ�:P�m}��A��⤧nJbR�Z�QFk�˻�RN�D\&OJ�]��`g�� h��-BŐV2�d��~?'��,R�?�rҩ��[׊��e��-�d�o��%��f��հ���̦i��c
�+CLsd)4��k@��6�u���s�PŐt{?�v'�36[\T��G���H�kR��B��n	e��SK[0T�v�d�d��N�kG�y�g_��暠�1&Fkb�A���H������W��&$�.G+���������շ�*��)��*�M#޼�i�ч;"�D�&>O6(����=�݈^z-�0م=�_��F��˔J/�����!���P�qo�T�/���$�`�L�Kz�u;/y��J3��Cֶ�&�3O���/����֨��A!`%X�jSj�'�\܌�O�Dﻋ��C�� 䟱٫��x�����D{�֠�|�� ��\=���e��G�T+�v�#��Es[{]s���"!F���
a�:�2��o��Ϋ�6�p�'\c����1 =��y{��_=#|�����?K�npN�;]����m����d���"�YA�B���n��n����u��]�Ғ�8]�F����K�h��<��&�3lG��ZYPr�T�둛��-`�U�O�p�܂߉V�C��Vm��9����L��D!��gXrA�bJ���̞!`��5��2�Q�_T����*�?��\m�"IQ����׹�c�_��������3����>Ý��E�؄i2;�d �$0�/��nj3�=�d?�H��[G2�H[nL0g\u�ϳ��z�%+�*<����G���V^�Ⱥegفt���7!�h�AT(K+ A�M���c+{���;���wa&~��9�/�b�	��$�A��F�a�x%l�|�B�g�U&��-�8kK�B�(��u�`kГl,B��q*T�3��2@�S�Uˏ���P�I�^h���RC��ti(�P��/��!WlcG�
� a���Pm����L�N��F��	��.���;�߲���6�4U-.'�����Y��m^ԧ�#[��d�H֙��u�k�+uV����u��=��,Q�O��ޒ�Ie�&�-b�S��f2�BY��D��.��n���n|ز�w{���j�:ާ������\a�i�*�A�w��i�?�쓙T��k����j6Vb=�Nv�i��5Z�Z������aMu��~�1a�䎥�-���7��ԓ4�Ľ���X��{��J �����������4!W���o}>����8�oɗ�d`�
�*�ՙaR�����+����;g�R�\C�쪵���S+c�Ѽ�>9�B�E����	�)�fL)����@�_k@����VM]#�{@oW	��p�$({����Lkn�>�.a��c��t$��c�J�u������+�n��a_-�Y��o�>����'W�s�B������J������s&���K)����Y:8HW�׃t��"���%x/|�y���������G��09��о�zӈ�*
�}���ѳ�B4ג�
qN���;i�	�,��m�I[��=ܶ��IWW�&0*x��+�7rL�����9̓�x�5�_4~�6b����f��gT_�P���)$���^!u���졣���޻v��=X��*=�	�����f<������v�5r�5ؓv4�9'd����|�:	��kN����H��ڝ�ߏ4���-2��S5$H��~љD�U&VN
J��#_9ǹ�'�R�
h��/١�3}��7j���`|\L�R_}�v�ZD��vd�p7�O�:�9�q�3}��
7�%"@�OҢ}�i�i�ǧւ��yg~������F"��2�I����H���E'�*�ț����#�dM鐁I�Pn��-�9L/ �>J����]Y�����������Q��%&q�j�X�8�Y����{���s'�B{���9��	���K!Qh��^	����'�7ʝ�x�pWt��\�6uI��U�[���<1�^�Z����W7��`%��A�������v��B�o���Lh�*5���m\�
?�$�oY�.����eR�[q���Ҹ��4s.׉�#>�@O���$ e���:��ֲ:�4Qq����v�5��uU�X�3��m����,
��
k0��F(��;�.&3Hг�#%ߥP��%ݩ�Z.��
V�S
?3����ݸ�W"�
�{
�[����M��G��8���񣻖3�Z��X����l�n����R^�<�t�RP�5<w��ˊ!�2�������;Q?N��@�� P(��1`���^�]#nY�$+�9�N�a�F�T]�YVz��Q�
ǐ�^"O�c8�v��r6�HcȎ+ =w�����#Ck��0�W�K$�x��6)c1����
��G��5��=}�CZ5��w�H�NtV/g��_��x1
�5����͞�~myu�1���o�Ud��%��1Wq��B���Vݾ�[��RB���z2���8�G{w���
3s��o)D��/��q�x������Ƀ�Db��ԁRc?S�a��@��A���n�p��mǻ����nf ��Mb�,)���6_��V�;t�*I��f�Xݧ։�Ǥ� 
]K�!Qt��t�A�W�xv>@S��Y�}�eb7�u�a��d,)����ϊ�%6Z�"���,���H���-A�b�yo~�9�ڝ��.�W�ee�����=͕�W�:+���F���_�%���v'��n0�#����#�:᠃gG���bD��t�B+uJ�j�q%�5��-�$ 3T,/Wҥ�^���O��W�d7���&ij.���1�G@'��w#)��sYS�K��P����0���!����I(����A�������Q�en��C%��h_�2u������A2�w|c)��
.A��E�"�� av�2)����Hi;o�S���4z���N�0I[y3y��|3�ѭ�+�O�
�#V��!��._��8�O��W��$��L���p�چi��h�
��5�X��[��z�U��u	a�Fp�0ْ�]�?/�'����a�ͨa#r�I0�nE�r"���#�G���FS,�*��'!i:N%5=-�>�*��`O�k6󯆥L(�)|����0=4��@�=��ٯ����<lm�`�V������Q��[r� �%Z�G�Cz}}�Sl���g=�,LTU���~����>�ۘ��BIL�A����U��& j*�ƴ�r�^���3�8����޷m�F���#.�O�Vޭ�I:��:g���~- �7#�U���?�Nê�l5��������<���z�I).�/���A�5�x�j�l���?�%��6�Lr��њ3ME8��~���V!%�#{�u���'N�EYN-km0����l�:��?�����/=J�׫�4}q�+DfUU�e^��Z�X���O��ߪ�]"�����H��3����]䞠N)��v��~��!Y����f���I���8��S6d�r�d��`<w��,!Q�^�M.D��a��k���Ak���	��o�&��]<G�m�RҊ����X���A�L·�x�g�;���&�T$8sN7��@mw���m�8�l�3JdY=2����L��o�e�&T�8��:�F��'c3�#N�*#D�H�X?�u:{CE���H4��d�;W���ǆL|�G�t�;'ľSh-�W!@�Y�Ed���1s?���Z�|������6]�1�g��C񦃤��
��@��6����}��<?�0�G���lZ�gO�\ɚ$tc�}��7��6�%�q�E�!�Z+���V�e��ߡ]���
���2E�L�w�.��
aG�~����mh�)��l������c�v�M�]*<\�4{n>��ah�@ψW��C�
��#��{���u%h	�ļ���9X����>���Sl�����^1�M�v>���k4)�9�j���g��$=���W���5(���|��xyDj�Q��5y�V��z����h��-���J��0��^�'�IU�t^�66�3�S���P~�yk��s��jȸYӛ��jq[%\
ǔQ��S�Ѳ���6��.�A��^!.$4B�-Ҹ�u,�l���>yS��?�[N���[D/b��,��*�&��z�*�$9�;m�`e&�x���&ƥ��v@EM�O�9s;��.�	�܋��� 'm�gJX=�pl����ע��ϝR��u���F�m�� ���+�=�%�BAC;�F���Q2 g�����-tyq0_��tT��!q�֖�j�3���G]��P:��&��W��~��pp�,0M�����4���"9���wд��}�"
W!�>7ԉa��t��{^=�� bAj��6��)߄5�apqߓ�I����O���ؒ��G��r6�͊��y;P����/N��`��S�Xw�Ui#B"\��.��>v��/����DP���t�VfL��CI�1m�~2U(�1�\�@wcC�=Z~e��\��f�u�¥g��N�V��^!�B��?�&��[`~7)��O3=̊�-��L��9t��RO��P}NV���%ͯl^�86�x������Q��?�'il`��@���i)Bnc���ߡ��Ah�~�:��KK��)��������$�*�j�?y��9����!�;J'��ԉ�%��u�c�_�y��?�V���c�����ǝ/�aE!���_��
��g*e�������Ɓ��@�=�]8X|�zY?�u#վ���9遢G�dvt�b����z�:f��}�B�9׎�W��n�"�`�ZUif�āx��'������'���IU��Ӳ3m��ϢV �d�8�*�����*�]#��D�����\�w #-'�����lmN4N���z��ܙ�O~&�x>�
�!�U!��	C#?�	�a8L�!���3"!/��#+
Ό�ܣ��*'d����tta*��S���V"�L;|�"B��v�*�	���j��'��
s��QzC�ꍑ��2�[j�h �HM�`�|�&�I�8��TwGY�t�A@`ְ���J�{���22�rŸ����W����������(8���ʧ��cւ��� �wP6hס��#R�N�q�����M`��"+O��i�}��2����6{t��;�G�9���h��#ӃlQ�R���m(�^�u8'��ʀ��UR��������R{�����/��|U���%m~�\��\�aފ�%i��{����H�ݜ迸9b�T�l\r���`��,C\���.��bB�T�n)�_!dz�c2�9��^�6*!��x�+�kД�S�X)��FA�kr��KMe̕�1�I:"jNK����"��A�,��]�?�^���D���b4����XqF
"���
R3Ʒsb"��ۚ(���} +��U�x�a���(.{�P� R"J��!s�KhZ_�7>!8QFt�";��8���܇�CQ�l�C�Z�B���dpv�T��b����V�o���,8�k���q����D-m�j�>n�����s�4���ǝjAؤ�ϥ�|��v�ߋi����0Y���d��ǡפc@@����s���_Y[:�/*���i���4���XL� ����'�����B����K�HZB>��T��.gc�J��A�>����-<|W��	�}
y���$KD����y�ǀy��O��T|��w�8'yq�<�go�h*��DYCH�F@d�I�{FO��3��`%A{��!m�Նr~�޵0aP�g�Wr�P�d:����N���<,��Oq3V�#�w�^�J�o�3����7U�+��*=�D9�5�s�j=�E�,���K�>�1=w]_F ʸ�'^��������ʺ9���P��2�4P� f��W��	_`�,��/��g��`��k÷���@��Y]�E��������)w,�)�XU�r��;� ���؍1��=���b�4�M��ɑ:�nǶ��K/2%AR$B��`2p�nc�O�*@�������Ͼ�C@��F2�d��
L�F+�i]�c�;��y��M��V��KV@Ͽ�ύ�8�`��v$�E�,7Z��$s�n�eo���n��ɩ�!��
�-ڋv#E�sk�q��n��8��1>�
���T|�X��B<�n��z�u�}�d�"�*]�E�p���ϭ�
�v/��'��0�Y_b-�T��]���+Ҷ��Ɨ�-�a�Q�i��`Ȍ���N���%��Xtvio�(�P���
�>�l�8�	����v�ע
Z_6t&1g�*��@wC��Z�Qٟ���:(\X���q1��"X��+��o�ࣼQ�'IL�m�E���Z�����t��L�i�U?ˆx�o76P�'�(N��W�~�r��[��@9\�I-Q�J�}52���awld,z$�1^c(;�ة�~$Θ�IF�&,���T��}��]	L��"}c�^_�ȸ{~�x%��qfW�w	N.�j ����l�g�9l,����D�]�b�v���6����H�٢�q,]���B2�����''#�H*��6��D��aŧ�W�<3ٮ��6��������]u�VZ�S:���LQ��C��>��#ٴ��%,��L8�H����X������N��"��}+4?�Dx6D�'_�4}#��?�/���y�࿥�.���s��kȉϙ�*��b�U�$i������H�V����1̽
�"7��X��&��)p��q }���棦E�&v�'�6M"5E�:TN�sZ�(V�=g�!&F�(0������Z�r����~pD���(*:���C+;C����i�"�����D����� ^�]�,ML�@���,g�"O���Ca%�A�I:`J��ߦ��p.�Kʥ�q��t~yG��Y��P�P����o7l ��
��K_Fʽ?���Z��^��_��
5�8�dۧ��A�#	�
�LL��H�W��]u+D�Q��a��DlʶA�0<CR~�y��n��ǕkS�߳cmIp2✯x׷R�U����}��
@�kHL��2�Ъmd���ʗyC�lI9��z͉����5`�����NDvt�����f�6[�b+s�GN��? �
[.Ȧ�.kJ��R�4��%��i���^KY]w���;MI?�}�|��A��8��k6�\$�N��6��n��a�X�:_E�g}���׻�iX��7=ޯ̵E"#���$�����H!���߁�6�[��՗"e��,���|c���I���Y��l4j�$�.�A���!�F�d}Z����Ynj���uz/w:L(��V�Z���}��^��Myr9��N��s`8a-�`=z�����Z�8p�ME�_���2<���MK���Vgm\����z��߿��͵�[�j���MO���i����U[���YxHm�v��4[��׬������-'�O��<H����e����D����,�ڎ�S!����Ve�ɯ��N��A�C� �uIY��ʢ}���ԓ���@iԀkwW��0GE����R~�g��')��h_vUp��Ƙ�k�s�J�-�7��Y�����$|�X�{é�����ߓP�Y���>"�%g�?-e��>͓{d�S�ޡ�t�P���l��(�-��v'��ù^��WW@^a˷Wa���0���zU��>�����%�,��L2?�	mdH��n��_G�5AD�)�z�bҴR7�fQ����G��$H�r���/�o ƾ�����[��xsR��ߴNbS�ȷ�}�|�O�#]�.k��h0!_:v+w�|�ת���3ң�M6).�]I��R "c���<FT�4��McUz#ϻ	ϳd_�I�
��y3H;�� ���<�Y�(ީ8v���=)���:fVp1FbA�7a#fHH2�_wY�Xl
��k|�E��{�����%��BY+�
���yә�{5�f2u�����B���MԹ}�b�;p�͉e�|~<�搒1c-H�u�C���*�cz���;X�T6`UEWd�!*g�����x�m�h(�XjHJ��Ǣ��[��&l��$� �j>:5�����>5�hc@����.;��_�	�4A'�%nt�qB[>JM�W��dz���T��
t���ZrG��')�;uJ��+X��	�c����'5���>��x�Rx]�lt��\�E�ʧdY�'AUb�O*4yю�,�nW�il]JS���B��N����ܰ�z�Պ2�0b9&� ��~8��c����\��J�s��l�V����b�RQ��ˣޥ&���`�^W�Z��/:�F��Ύ>�@X5���ݼ�9���O̩����S���\%b�#�q�uF^���%�{��ףmɝ��?�zL׽4ܞ�Q)f�4�Z�{l�(Zܖ� q��[�z�K&;\]����]/��O��xB�<p��2^�Ϊ=�{Q��ZI8�$����a���z5�$q��+��#�����c�364���6�+�w.�r5Y�[a�Kj��7���?�-k�������l��^�j����>R��D�~�k�>F� �h�Tc܈�$��`{�',� ?�>p�${�A+����k,��P���{iM�dZ��ܙ͖���0�C���!�:��Ip9aALȭ=��oΑf1g1�9`�&;J`W�����"�A@o:�΁ ��%���d'�HӘc�V9M���i.���u��������������S�����˒egɩ�[&������k�p�	��MT��m
B�����/	�����|W`���k����Pź��XNc�&���k��c^o�����+��2!��ϔ�F��i�V�;�6��*�"��d�|��xy1��3��1���!�y��*�8ť�,�rm�	�Z�*Z�	܎���>�:����MTk�@��Wtn�Jp;�E����c��K%�3����䊓qRw}��f͵M:�|o��*��ίH��O��kp���Vv��25$7i�ZN7�k��^0iD�o�%P�dke�2BGM�"�Q`�?`�����H𡍍�����Y9_w�眦f����3��B+��ˈu���֒ɺ7������c��o3�U��&Ş+����F7d��Y+��t���6�!�<���w[q���G����Lm	M]v�����,��c���S�X*|���z� ��a9�,�k�|U;vK�Y��D��P6D�@�|:]"��MKKxѶ��4Ov�?�. ��-<phL���S�,IC�/��e�����۶E�'*]��ZVwS�"�$�����'�e�G����t��RR�`kb`?\��OB�ͅ��ƍ4��z��x��7�4d�e�����ͳ{�:��1���^��h��n:��i5dMr����YSsl�*ͣ��l��R��������>�Bj��Qp�1�=��3�]+$^i��L�%��*7�c���,�Y�!I<T$�j<~��@:Sj:�P:�§�̩%�`�4u��V,)�H�A�l�"�Ƅ�M��2]���ryR�Zl���웎���βB�q\SS�y���2��0���FQT z��P&w�9�,Ҿ����8@aZ�\r�;�4��H10�y�&���2��U<��~�����]��+� ���O��vh�R�w/��h7��sEj����d�僧��Q�韙����8��>�q9�;;�#�uvi��v"�]8�>eEA�5�bi����/WM+YL�;a�8`�)q*5ԥ��4�������B�"��2�ۈƉ�:E�=b̛ψWٳ�r-�8�X�p����T��R<��!*RX�̂�K����~΢y���2�v��۾HB;�,U��s8��
��=�{�O8 ����`��uF��1��/���v��㣟Ǯ��\m�R�a�=A"k��7�8s����a�0��.7s/�U`y]�S�mr-�p;��m۳�R���H��K����v�y�A�����$Y1A$����V����!}=
vYX�j�Օ��s6��L��f��x_	��c�3���\c�Q����|�%"﹧���ʢ��W�$�6��	��l�����]���(��CV8��������,
��w���p�=�Jgz��k��j}�e�Ĝ�+��AY���v�;q4����tN�4��fșiݍ�~���ސ.i[�:kA���?����*n�2)Fu���+b�B} }� Q�r�ւw��f�'A���v 4֮3Ͳ��1b�e����T�WO��=��� ��_[�\O̰KI�yr�s�uɶ ��/OXn���+��AT:~^W1�=~�Jv�[�(.��F�D�H�p%���7�KԖ��}?�����E\Z�����CV�?Ey�� :�5Q��z�&{��\b�K��yo�ľ�a��,:���Z'4�uPv����i�l3J������v��rw�"��nC��.D���V��^�Ǐ_{N�x����D����#�5��b,�e��^�W�B[��81�v`5�O���q����@��@h��Xr��Qoe(�50��aۋ󲆩k�)4Ї�~�����R[n�m���z���6�7?��ߩ:�����9+�]���%��T폞�\V�L�̡n��EwnFgt2�8(10ᰦTX���f/�E#��d��c��d�'`R�F�]�qw�`S���0�"�e���O�"��oz1���=\-ҋuD�շ9��̠�[)��A������DͿ@�*���i,�gޒׇ�l�&.q���Yz܆�;��h��U���P���矏�y�m����-�r8��&�G�|����@�ЇH>��m[dD�^u9�=l\S�#V.�ud���u`:͡��6O��)��wʓ�)l�Nw"\���Ɩ��n�~���'i7�L�*O�Bt��w3��#�h :��G� m��A@�j[�3�R�ͬ(��6P���.�L��CQY�ͺ�"�4L�s�W�q���d܅۬%}��M�j��˂_���X���ݶ��|�d��w��q�Oe����;J��Dm=1�s>Q�F��)	#���&
?�2�'}�Vu���_Bn�������b5w$��}�����$:,�4�yw��`�ĥN�Ծ�&���΀�mߧY����u�ks���^_fG�nt���~�Gq�sj� 2�c�4I���;&Y��{ex�S���Ƞֶ��}�"��nHRra�8��9o��gkϴHW�/�Ei�5��C ��<0h�N�]kO�x��	���o����=������|*���̊!r,����Yx�
�lo�	�|�C{���=��8sD��,��M�C��j�eb=%e!�����c������2�����:D-�����$\�O��oX�{��!w��)�@�{C�/0���~�'F�P���%K̵{���s��_�MО&������)r����Py,)+D�|�Sl���ԥ�v�V6|���llikO�En��Aq?����x�`�K�&�7�0���6~@�|Uo�f�����~��p�y���F8�����d��<�M�>*!�z���B0�ΣH����jHIF|5��O�b4_2 �G�b�uq+\�\�0 ���=j�~T���q�C�Ѝ�����p*ˀ#���V��6�D9�>��+s0��?�R�h
�y������<�,޼c}H��,?����{ k6d��d��17=�^�����2���:�59��2U�q�	 �)b7m'?�̇��xRNZ3��qk�B�ʬH��i#��m8�4>V���Q�Ǖ��r����;� '�r�Nj�J��Xx���CD���zwP�.w�KD��]:�S<��s�S{V�������W���H�md��F �,g�{��K����;�Ks��jy��M��r֎}`1[����~\�.Ø�yg9���b���h�6CK�#3����R�a������c�}>v��i�K��~�c"1�V=�bA3�-&��΢JT�!��$q�mb���/��H�C��W�?AI�M��}C'ɱ^�hh]���3HF���`�U�7sq��X���ؔ�\�y΢)�|q�>��}�#W	~;^/��:��B�T�3c����޸���x�ԠN�� �8���\�%'��d��������d�_EC��[�p��b�>}���8Qv��Fx,�<&����>��ù5wJ�*V3�/����[�;����e暁`����^���1���{w�yJ��3�l�Ba2�AIp���_�cR�y��!kL��TzV��D�߁�ݍe��YY����$�z�%�	�F��_ߞ�&<ur)��,#��I���S�$�������O��	�fT�(r?I��`�p�
l�i�|��fb���*��R�O �0,ds��[$PC����+J���@�cy�H��A�X^f�����W��bD�/��C>[F��h�`)�H� $�����́�5�kVҪ�Q���B��V����L�_���8�����;�|�^�R|yҾ����sC����q6v_ik���E~��: ��F����<�����9_Lt����:�o5�:�(
fM
���,9=1�����
�cdDCh���K���Z��jO'4Ў B�� A�3���K�e�c/��ym�k�
=��#fw������ ���j�UW!�^�H܄�'�yn���ýQ�0���V�nE��ۂ����l�	b1�pױ(j�H���3cB\�N?{ޅ�:�+�
ږ��UKRH�8��V�zz�d��'��F�кQ�!������5c�&#�la%/���u@��r�v����&̒ :WLw�͚=�<=��@�TSz�~�F��wI9��[/zN�?�q/��o���)?" �Gl8B�����Y�eK��y0��戚B^�t=�P�!ʁ��O�������"��/��L����m�ĤQ�_���Քt���6�<��u{?��d�b�u��J�	�>ܘ�]��H}%G ݄P��m��/l���key���M�Qp%.i/�̸8(>����e���!�߃�q������)y��!^G
C� i2������c�"�B�ȕќP�Wd��vmH����T�C%TJZ3͙���:L�_l����bS�xLχ�n3�����{��H@J-`[�U|oa*�OHZ�Δ�=�?�O&��`P���
?*D�7����񟄞˟��u��
��tSeҿwRզv?�d�xS�!x6��+𬦜x��Wm�D��2��~Г�qb��8�4Д�Z"^u��ι��X�]0s��T��m�o��k�W��/��b��=���$��S��y܊��	D���ؤ>.�X_jw�&X@r�7��2���� 4�2\`s�S�b���c��{B~�KҨ8ݎw��}%\1��nՓm�'�@:��m*��Z�+]�l�eg2��E��[�z)��s_�-�Y] 3F�z��#��/�jf,@�
X�eJ�u�|:f,:(�S��κ6&�]�3�M=@5VN��%���G�Wb:m�{�Y��bWNB��l.���=��f������7jwroA�JP�����@�����s:�
�:��Ә�#&1e��+S��>ɞ�������@�N8r���عF�����z��WW��ϋ���T��F; || P5��0�ʅ}QO���͒I��a3� sOk�ӈJ-����,�>E�1�<�^	�2�Olz�)����E^I1ZGb�C�6�њ�c蹱�$�^�����ܫ�[�<�h�q3����py�hY�p�'c���x�Ӝ�7��P- <n7:�Wσ��v�F#\N�fJ������J�}�U�/��Vd�>�}j�ӣ�<'��e�r�}�9��W�zC {,[�GW:�m��35+�����%9-N��.��3��k�Y�Uɮ�<}�8��q��v��8�1�<��#�)=N�Br��F �S]3�5���G/�N~7�by���{��#��0#x��j�'9g�C���+�����g� �J>��w>K[8q�VMu��\��*ZQ�-I���*�E���Cq��y
��aK���� �fn�HcIz��o������+�=���$mI>�8�G>�ʢS�7Nץ�/b����-��.���ZH��&��7¢�n�h5�D�z�t��_�t�F^��D�B2� K^}]L|K\�|�}ơk�wsu�@�hF" Xp%I�h�z��A��Ϊ�~�<�vG��_a9�<�[d,ee�f��}�f��0cyU���d,�n��؂xǃ펶��ӰOTqJ�j�A�-h_٩�؂z(&���h��-�DO z�gv47�[�>^�ۣ����Ci"��r��`��_�g�Z��0p���>�FC�������u���@�����"�n,��K�6�K��e
�����YV�:��Y�/'ӎ��U��l��At(.�!A��G1�)"a���Q˽x�E��J�����#j���QL�0v�MbhZP����X��0������Z�ge�X ��Ub�+(��>)��Ƨ^Pܞ[T���l��\�e��(g�9.�.]*�3�����N�Wc�âs����˒3[�_{��C�kr2�lb9dWP�|�����!��d
2��X�v!���9R��Y�n?� }�n�X�D���G�U����}f��'�%0Y�4Y�:��tn��̋2�"0Ĕ���q!��Z}�:�C��~K`�uo�(������|�cR��yɼn�� b��	~5��R4�`J���{��i�q
�,�� !<u�A�c���"���	�4ă�ẳ_P��ÍD_��-��#����.')��j.9���F�%�d���cl�&X�A��2J�>���q�R����מN��c�3�u�p��\a��� _9({�n���U�L�7���ߒW�J��\!n�$����t97�ߵ�MU�ne��#�`?��YܮI�9��^;ov`q���H����;5���S#8@ ��t��.'��$f����S~zkk��q�<HI[Y�t �ɧ��}��A���r5�?��VHĒ��v2[�7S/U�m��S.���/?5q�P��X9�D�w3�p/,B�+�	��ҋ��6.Шrߴ��`�~KCυ���5�Т��uۘ�?X0]5AR��^TG��4��gx`�"��~�ܢ�_���w�@���lL�h�K4�6�/�����
N����G�o	e��t����� ����eT�U����uǪz�=�	��Y(��4R�3çH,sYu������4��X���}tM��W`��xU�W����s���c��zx�/#.����:�����1bt�WS���m�-�Y�->�H{5�<\�:8���}�gC�)�6����$;���/eM���#4]�bP]r�j2Ƶ�༜l���.}!�Id,��2��>q����Ԋ��5mSd��d�&�,����(�:x�L�Ò���Xu�r���-8�o\1�o\rt�mbؤKVz��у�佖W��/��*�_n	ٔ����1�1�6�W��!w���|���TSE��.#���`s��*�9���O-��D��2�����:G/ׄ��wIq�0����y|���͞�| ��<X���{z�un*�U��&���	5�-���V��4	kއ7c�EDF���U�;����=��)�����F�(����IkC4��z�l�$�n���}�J���Ou0�Z�f����
��x_�[g<�hѕ�����:ld	���H@Y�dH9��lsd����a!8Q�$�ِNq�G���@���-fH*F��|���,����Pܖ$�3���ΧQ�<�pZjؼ�O�Z�ixT7�0��,:.
�;�;���� �WP�����C��`X�H�j��N�Λo�.2-1�W�鵤	����
�qi�Ȼ~�o�S����)�A�rO�R�ė�hI!yI�$Q�K�o�������ɤ�9�#)|�#���D�* ����#����eI]#����S�}do�z�wda��B�7q��+����k$V��J�y4A����N��@��Z�`a�}W�� g����!q�&���AmP�"�]>$m�
�$[����� f{�O���;�C}�T �ʃ�#���΄���.���	SA
4��xbd2-Q�	�el5���=��2	<j���vC��E�v������=����3G3x�+L��uu0m�rC��v���FP ��Cy��O�$q�RfG��ǑV�8a�X��Ð�.w�G��y��&L�g%�4�v{�\��H���9��gz����%��2TT���$������kR��T��3�n�����V������:�/r��|3&[b���Ĉ䯄/9T�ag$Ӑ9VjB�JxMzٯ~�	8�y�`ǞO`=*�>!c?��F{�.�k2s8�`��(+����*�>$����Yx�6X� �>�y1�HE���3ڒ#L���-�o֭�L�X=F��Q�Ӻ��42��F'���Y���`�*�ֻ��2������^���-9�8��[pH�����Ǉ�,��q�%[�t�O l��9")eg̣��HY�b���
Dt��8s��)���:J��_�Ȁ���,e��b�v�9c���m'�A�B �q"����0h�7������
� � �(�C�[Q=�M����V�jz�����>�GO/����X���m'$�A����28v��G
�si��yYǺ�LT��3�b��*�Pb�"�?�rцQ��w��)�е��MÄN�$,}J@s������F@�b����y�H�$\;{9��)��(88n:���ώ��_B�m��d��X��%��u�L��ʢɒ�=��s��������Iq��iP�B��GƃlG+9;n�nM�r�|����Y_����r-����j�8�5�H� ��V�@�x��<Ѥ{2�Q������ÎX�K��53���{�b�ngkޣѩm��3��&%I�Oe/+��6L2�.�+�r'춢g�MjV#T�3�!k����$��!�і"�GB3��̗�)���z����~+��*i��}7T��H2i��ۣ�#b��O7��A�$��qL��ֺPd)���`� �VU��h�Lj�Z�v/e<e�|�b�B�#�rz���h��mX��	�vTt��8����L�с[j%D `�|�!%AV���:`焙U���Ā�ZU��V�Z���#�O��2�D�/#%f�D4m��3w���,�K�L�����Q S__JD��f~�ܜ�r��@�=�A�Մa��`\�o��5ʛ�P�I�$'Z{YJ��/B�DG
ILot��XѨ���ߞ�)�KЬ�p@n�cj��ڦI[_:��^�ĦA�Y��RPk98F�I}/�yq����k(�K�i�p˳�3�C�MM����_��d��O~�뤵s.��4�P���C�����旋�/�U�o�e��J�����Z�csk4�6��Z(hQ�l!�)Eg�DL�Gu/�+����SD���_��erU���J�2���?���{u��]����,�����/pZq�s9���~��s��%Y�Y�G�hK�&�N�Kr�]P_%/�2��j2S����vݎ�aGq֮���Thc�sM&ó�ert��f�=�,�A��|��:^�4G�XOF�qHd�>�؉��fdY:o%��%��X����`yF_��mha��[�qEJ}JS��~�#�o�P���r�>�j�P���	����+�+� ��k���0�[a�6��7�=��� ����0(��3�wy�
�v��`Գ�]�ܞ��h齡���.�a�RMB�\q�������8Ѣ���:ΰ�P	e��f�	��'��0�Z0�����d��7�f�'�hE��#�Kmm����灶�+h���9�͡,L}�~(��D˸�֔	m��pIE�G���9��S%Qo���K�� �NE�VVɇ=�%J����T�!c��Y�Kd"Òm6�E��!���vt��n>��?*pz���CڭSҔ��U~n�zL�9a_6��aH�$�`7k��NP���Y����Y�������G�|���f6��;�ʛ:fͤ�Z�1g�yA
�m~��	HK%�]�����=���n�k��J6�b���ySe
v2�E��N��&c��I�upDy�w�L��k��Xg���'��@W�~oq�34!Yݸ	�R����6'*R�$u=#�F��#�;�J��k���"y�x%�:@v���k*�F1��g����o���q��=��{/��g��+�i�Fnz�Mv�O�t��>N=/n���W��&�9���A� 5<��0�(6:�R�)�7��4����Z��9v)�+��c��'jtLϠ��F�7h��!��+��o"f�V�+��u�!��؝	;���*9���Ϛ1��n�E�^�Ɍ�UP�d�7��/}Mp�����x0�����V���j���ׇ5�i	��3Ms������U�¨K;Y��b�p���~\z��i�g��R�-�/ �0�o0�m
o��࿯Mv|�6�D�j��M��u�AU�|��"
0�oC��O�s;X^1^���֦�LXN�
�V��a�q���/�KR0�i�.(��1��Qu!�/뤍w/��qs�+R0�jki;���ں+�ϓ�b��:�{@�ܵ+Ƌ���О�#� )�� �3L�S�J~&{~��9�(��G�e{�߰R�s�iT���ّf��V�����3��&ݭ%��%Od�~�i�s�:6eK��^}ή|�bst�hv����������ְ���?�cϚ�桛��| ��
����f���	�<�,�t�!\ E�%\D?(�7�V��ݾ��c�1���6V�Y�M.�$���������8��k�m�+n'K^���/�\���ց%iS,gV=�5�	xl� X#���MxM@��i*���3ޒ~�"{ �E������lY����5҈��=J�,QmA�mtt�UX8إ�6�D��N��fk��A?%�D� ��p��}��1��1"y����ψ�mã�q�߸p�X����Um���=�>[>-4��P����ԟ�Hvk`5��^a�����Ϟq�qL�O:�7f#����F���I=ռT����]T��0����PO�BO�X���.�N�C����2HA�e�:��o�1^����=��sU�[Q���}�ht۫	F�84��6}�5!���$�8z[��8����MiC�H_v�f>C�V��Q,A� ������Rn���Ԃ�{�Ԛ���S����ǼA�k߀g/��J�Qxo�$7Mh�|r��$7�������O�+#�y0�-��KC�� -^i�l#�����_�Y�P��J�)zb��脑��������Ã�׶�<euVȤ����� ��g}�Y��R\MD����&��D{=�������]Җ�.}���Ry��똭=5��!pʮ�}��iU��A��7����["�=,Q6��}�2's�g�2j�n����D�^&��Ly�97����qh��~R!H9��gG79�)�`�Hl�Z�8�H�PV"��z�[�G7_��	�㺓��$�����-���2�s�E�Jn̰uF��>&}��;;�W x� Y�0k���A&	_�1� :�f&�ر�Ip��.�����K���&v���#diS��nI��K�z����1ʈZc&y��e�n��*����ȷ��š�G?Ƥ��;�%eXܖ�LdQ��(��?����y���"ڈ��9S_4�R_���*H.��|T/@a$0J9��R�QX/���GT��G9���]pEu���Ј��g�`����7�~���hC�%1+6w�?���^��W���u��W,YC(��u����i}f+�b�Uw�p���y
o�ƌ�Ɲ��<.�.��dӔv uh2$X��vՂ;�A%q����ڽ`�>0�G��!5Y%	u(H ��������r���߀%����e5�r>rɏ8mTQB�?�BmU�`S�Is��n��8��s�����[���� ��o��O��ƚ&4�6����+]��Ҫ<(	M��b�1������7Ć�f`sq'��a��ėC���#��@��f�1/��ċ��k^&p�tH�dy����Zp"�LƸJ�E��06�}Ҕ�UZ����Ҿq�H3ΰWZ0�ىPm�ͦ;~kg���$�Jt�re���!�k��'��G��8���?�i/��3W��2hκMn>G�h/mP��IM��y�L^����מCa 'Z㱪�X����J1�^�ܚr�������:e�MI)dg/�j��x�o)k������7�p��bBeՋ�~�+��"���>��^lt���]�}0ϱ!jlD��|i���}��Rڶx����O�1|�p[a��K3u��Uvx-\��*�'8gPCy��U�nQ��|�����]�А1��kcrȮ=��3ʯ�Bfѧ��Zl?�I�?�렢v�I+'!,�e��?��o���Vxy�9�N=m�q�fd#o��������i_(�'�RT�]��U�1���2ȇqp�<�E�ȍl����.��VF�_ϸ(�w_�nԙ��������hLF��_��l��޶^.��6桺��@9X�ļMy�L*e��FII��3�z��E�|A�Bi�l�:3� ������%�+�;����+]�J-t�؉��;��h+���]��H|��^�.��QL�BJ:�]Gye(�m�.D�{	�ee�g���/��S��]AV6���'X��IuO��]�/,k���hu�xh͗Bӥk&cG�B��_Z�Ҡ����� B��ھ�������s��Ԕ�3MN]����B}D���!��%���&���+e?�X_Y�f�CkD�آ���� 0de��q�f���=i��k�����:z�P����7��t�>��48H�9�W�{r6��a�+���5�,���i�/��Pdq�,P'�P*��?�:��(0�[6VP��I)�S	�@��ǭ-��.
�v�?j(���B ն�o}��x@����
2��E�¡�
�a��եz�z�g�6I�P����QŠ��x h;�V��0p�lE:,{Ld����h*
I�e(��g�>�����c�E?F�e�;:�z|L�]/��3�\Lo6?Q��Y�_�D�T�!`�֦�x�I���Fs��T<�`���i=�g��q�z�������o�ͷ5Z%��9��&e��2�A��b^���2P+����0g ��=�_���[��lPh����,��{dS��]�G��2,��@q+r0��M;�|��Qn�0�b�1
.C��)Wl�`xĀ�L����Pl$|�����,�p����i	�f��/�C�y����n��ѝ}��6^_vw3�̝�!�ǭN�C�wz5��� �O흏=����2��q�:�D�o�ΪӮ,�#aϪ��c���>Kfx@|OĶ�S|j��>o�w"7m|\.ا��.q�O��2�4�,�.4��
��\�k�����uڍΌ���C�3��` \��F�fEv9�.�e��v�rF�Ù��M0�F��3�&���� ��:�K�;����9)�yTRR��,����ˑ��Za�"��m�ضZ�NI���P�\2$�ݮf��,���T���X��2���QNE1h����ENa�)��@��T������ �wA}D����%�E�l�=l}�p����Ă���i���N��-c��[�S����A������g�?��yF>�|���c<(�&��R�������[ښ�N�\w�p� ��
��x�҄����踘Ñ�0@]DۨO�D��|���� M����м�Z���d�̌��5w�d�A�U%&�v��(�����闷�!�z��1'ō%䥑
*��o$'A���������z�m�c �to�+t��ݛ[��<�}�|m�s
�ȰUC��[G\��Vr������k .�eG��	���2C;*�O+*p$mD�r���O'���0���#B
�s!�Z�zXF�T�i�Y�:�m��U	S� sيq�L���(C��<�Ȅ4�C��b,�Oŝ�̶��#3���l�������m5��9�f/;�4��J�����f*9Ցl�� ��ڜ�o�	�,�_�	�U�ҿ��2=�(���?n0ly���A�0�[l�\���y̠��^�C��{�C���I��~	w=���x%��$+�|�A�*�z�*mD�9���+f���z��^�U�'t	*!�r�ZP2:��.sc$z��np�j}F�ox�y���G65Lz}ۋ��O�d��^N|V�b��@;��2���n3c��\}��d4�(k���=>��(FAi���PDܩ�X�N)��O%������r�/����o$��'��}�¤�^oEF�4hz�]�Y�+%�q���U](*M�q"�B��
O�p�K[�M���.zJ���ĳEβmG��	��-_�r��8�*�*M��[ˋ�e�]���;&$�Cb�+쟲D��n����0�:������w��2xe��@� ���a�<��ѝX���sv+l�ixl��h������m��I�)�X����p�W�|�6��\����;b��O�֣�aI�iw�u��il��w�k��@���@�����ہj]}���2���50�E�F�~�`e^d{��l�L��N�N�{�u5���p�_ϋ���) ��h{}+k��3b��}Ni�̺n ��Ms��rb֓��_ eLc�]����稜��V�dW�Ɣ�ۙL!\��K���_��G��|�=9��}��t��`θv��{�z��c�'Z?�pjU��f�<n48����pr��Dړ]x�ao��!qLeȗ��/��@T�q2����Gu�O�����P�˵F���%SzIt��� R���_�f�)���P
�����9H�����)��|o<'.��z���N��|t$���@����\
�����a-��E
pd��Э��x���-�M����T�V/@TD՘��sy�\U��ߖ��G��1��Jg`k��3h ��&�\@�I����T[FCP����V-g��O%l��+x9��{�hzE/�B�-�VN�)(s���VY��O�tלu�A��s�˻��h��:CDQh��g�2����Uq��z`�`
S��=��7zV �_��BwE��l�|%��Ū�r��d4C�};�E!40�ЗQ�<�=�Qn���yܛ����������������绊ק����ݱm���.e�芙�|gL�"�u�մ��Ί�9�����:�)�SQ4�LuD�Sk�z�o�섨�v����e^�]��F��7.���ӂ���0R�&��k�&���~�V�X�k.+N|���5?W� 4-��9h
����������1m�.o�����4��[��FCy�p�@�iN����{c��%J�%,=�,�Q�b^حGa�t3�T��*�,с�`D,]߅9��HX�fxQ��y�e{.�q��%\T�`�A���_C^t����x$�EB{�Df���D����2�)҉C�l��r�~�a���{�3�{����bY ;�5���\Q��y�ruՓ̑���ڶ4���X��i�É�%�s �Aw�~+Q�0:
��#� ���
8�U��r�����`����8z�L�["@LgW��s��	�cIm}�P�~�Y'��4~wy;.\f��0
6��Ԝ��iڱ��k0Ǐ��\�t�7v���m~�����/��s�l��I�6��"2ʪ|%ψ�RoDE��Lp\#��lJo��I$�U����D���4H_i'j �s�i��\�����.C2�Ѯ5ܕ�D�A��r���DF�{w��Z�ԕ�Ӗ"�nRwṛ�C$���ӑ����".��C�'Ӡ�Ҁ"�x�?����~��?�9���6EN&[��8G��D�Rx9/�1��A�R�׉.��l�!o ����A�7�U~Cb�A�E_ 6q�J�^	��t�б��5H�ʱ�6k����`=�\�}�fǢG�X�R��j�:|ʞ�xLT(�k�~�!W��A;vl�|���^0#�����w����2�u$l�r?���P�����iݏ�Q6r����v-'���3�heC��k��i8��	3��HJQEA��B�� ��ۤ�@N��Ij����K��T�U��Ҁ��C�-�1)��L���b���l�3J��32odd����w��k�ʺU.���6�neK<?K&e�ڢi�(EQP��qR��~3�E�2�dc��կ���{�M�>����<[{m��<����n�P;����vޕ�z�L��N��u6����j��۠����b�c#GB�bѕF�U|���c��!�W]��ha��c�9�h�J-�%I� 2֊.���Wg<?Ħ(��ť�)_"�����_���P�����sGq�D>ƚ�����淒�
F�3:=y����ٮn��{����zdU��n�����V��K�;�O`�2T�2�*x�1F�P罭�ŉ�}�Zƹ�����7y�Ǩ�k��:'����x��\�#.�� /�Yå˸qX�͑��.�[�����Γ�ٌ��#�ã����-�^���3�
�'�t9�F��[|QSf-)ê�;�<�t~��b��oJ��3ǨZ��"qD��ʊ!?�-�cM�
�	�ZE�>�ZPs�܀�Rp�LY�7���t�O�y���~��~Yi�$�oچ��
?~Jx��ĝ�y��ׅ�XJ����~hu:�x]�%䎎z�h i��ԅ����x�u�LԬ5�R~�֓������"L�at�E��h
�x/<wxj���=�?]��.'pXo���Z��8ʃW�Ѻa��O��1M⡆�v���~?��6H����g��%�ث�����3��U>G"��XΗ�&��(u�p氚T�,�-�a��qCN8�.y��yD��?r�+�H�>��!z��}����|�����"j������NI����W�O�V:'��+ ����\������JkJ�)T/��0��Y�,+�5S3#��ە1���A�#Ӫ6�h�(��D�K��Jmv���߰g=P�Xjn`�!$��KI�KY���a�/�V���pM�өϐ?C�V6��#Oˉi�y������.'Ó�;�|�k�q�Pz��%�T�T/^�ɘI&?/��a����-eq��j��#�h�l6�C% �Ji�����$�
'�������:2#�͖�0��_�J�c>D+�e��\-�ŀ�E+J$��|�҈��u^1���g���AjU���q�6��W4�i_k"��m͍q�)�'BzW�h*O���I�و�MN�T-�ᆋU5�=;��B[Y :%�o���UՉ������!�'��R)�v9.d�|���f*b(�Z�C�j��ĶRF�f�r�����*�t潠�e"�..�g^��+�nIZ�j)Μ;*S�HZ]�X�0�5 +<�}4cg,�-�E�I����t<D�j���nGXf���Q��[���N�#׌����"Zb��cv�*A���h��G�C9N߸�
)��;���Ɠ�g6��"���i7�ST�p�}w�� 
�Y٘�Ôڨ���tV$�k�S	^�p��4Ȉ�
].)/��K�"�\�O�9����4'�DR7�M����l)�B���0!P|1-�.%�\Q�J��ge���ܸ����#ۖV��/���R��y�"L�/a���dʀ����	��ƻ����UϨj�� 8���A��E�+��?��7����d�Y����t�4
�Mfl�_㋦M��5���~Λ 4d�O,�K��~�**8�O�`kx�����}��!��sHur��`�f��n�%>����}�CW��HJҩ3))��>z�y	4����v������|�p*wz�A��g�n�g��a�XW�C͑���%����	A�PFZR�����{ o��]��|� ���[б�n?��l�T9�-_�[Ð�Y�j��q�L{GCؘ7���=�?)Q0	�SR��"I܂�U���G��8��P�Dj/*e��:�d��;�^���aş:6�0ȵ�=��b�/�����Ŕ)>o�d5>^�*|6w/#
�����w���X*�A�Bi���+.�Ȫ\�S�$�s���)����SHQu���v�-E�L���Br='�a�\�L���f�C��q3kBI����Ɲ����S���&.b��i�Z�;5LΖ���n������"�������;#G ��}��O2����]"�o2M�L�����p?��3�X��z���ܗ��� �!���,�x-�W�i����h_
7#z^���IX[��)DxD�)J��bBP ����70D���3��*�g��6�/��wL�Wå�+@���=���m�m��*��8(0�>v޾��z�/�MF��=S����'U8\����vw���h��6�N��MapO�u���F���Px���B��a����Y|��騋z~���v��)Ĳ��ޞgRSod/��*���h��]�?��lI�cQ\'�yZ:L}P��7�����a��7���O��w�����l��Qu�[���E�wSnfR��`G��A/h��Z,��ҦOL�a
�9�߿=Xc�R�j#�����U�9�S�4��"\�z��x��DoJ*�l���s��m
�>���%��lz�ֽ?������L�j����[�f��7 {�(\��0+[X���������A۬���iC��|UV�.܅���kǚ-+!�M� ߭7����u^%ޥ��@�q�z�s��p��"�6��:'ީ��M�Ǯ�U�"у�ϯPۊw_��Q��⢡�_���WF�Nc)�Ҝ���/i4@V� �UT�9�<�l�C��PI���n:dC6ap��G�霭���K�)]��t�Xm��6,�(	T���-6eR������~�&�=�����Bm`�3�#��	�?ʦ���ic�s�:҇T�"Ñ��oW���'U3��=T��IH�H�]�Zt���;�2����90Ǹ��)^\	t���r�՛Oj&*�?V?����:n�nXiO}��ʑ���lMg)�iH{� ����[o��3����mX%މɚ���C"�r4���o��4�S��J �Gd��zdSy������M�����q1���г����'ȱ���o��ӔA�뽧��:���X��B�&�rO��z��\J�5Q!~n.�I�Z4eBK�oA�?�?���t��E��}�P�������G����3�>����r��:>f9(S���m��R��W��K�&s����#�%���{�0�E-)�����:��&�_��[�@46��$�쌓��u+��Jd��?ߔ�9{���h���܄f�!���qlo�t��iM<����eI�^�*l�g�q�7���$�X�����ו��>�������ģq`��p�G�0��䁜^�~�P.KO�)��Q� �5S�������_(`I�d#8
taz=i�9C����~EV��	�����4�ܢ���Hz����y�%���?Y�"�3�>����E��s�(A�k�Z�6���f䬫�՜��U�s�d	�U}��M8��x�I���u`�2ssl��u�B�o.�V+�����WU"����* �&bk� '���z2���/U��n��W�pa�� ?�?-��1|�� d�U���i]=#��tbO���}�x�q;���t�D�A�ѣ��>��&Y;?X��g����$&�!#� ���t?�a����,Yddx*����w�3�/%/����W�!]&�Ͻ�U��.à�[L�>�>��� q�GJ{������@QA�b��]�E��bG����'�`���$��~�O�8�Uݼ:;!��3lj[�}�6�����߯kZ���z�#�*��o��QW�R0Ҡ-�
>��8Ot��e�M�m��r��+#�OR8�L~�o��3��s�'�����"Ʃ������
�6��|�!���WHW]��J�&9��F�d�`�r���vh��%I�,�ɳP�*�[F�!h�#��M�5��E?��A���dN�Zji����!��v-�H�}��Ixڦ�,�SO��W1I��_��m��2��AT��gR���"0P"o�G��i,?���ɍRiwɗ���&dA�ة�t�R@��xD���hm!/ߕ#�9��/R�ZG�Sb��M�8-��k�Spb����w��!�����@2"DNp�]���^�i����ܦ>"]*Z�,@U�o+�nش{�ە�cW��?�Ųq�A�QW^��?6�J"Gԩ�_Da�U������7J۽��rr��dS\�Wp-i��B��kߎA�����lM�O��1�O鿋A0���B&ȕ�,�l:�v��:a�p�"��s��t�yid��W����!��URhH�:��m��|ש�	��Y���!}�+M�0��*�Ŀ%��C���-�}�ǧ�Xn��t�9)���QX����|���n_I���G�J��d	����Ώ�b��z�4:Kp>��fQ�r�X��'k�{���+P�߅x[��v����}B�1�}��`QpO4]lQ������ӆFٸ`O�\_ޓ�WMi��׵¯{&�br��xrn�ujџB�^�C7�tx����-��B{τop�p����)߆FbM�7�cH>���:�����T�o� �{R�f�s:S��i,���!��[���*�.c��2l7K��04((z���oD����&G�}l�{-��PM����tH�UDjE�F�m�c9Ytk/��iƐ�Q��A=E�!��M9w�c�U��䫲��=b�M����/�}��ו*Nx_�ޗ^q�~K(JD��K�5�(�`�r^���	����8Ҷq1�)~"'"�ă�*�1�gg[`�|
u?P�\��d�qQ�. �.s�f�^zKgJ=g(���PqTw�yD�L�v��J�[9��c�El�����%M#w2A��䞡.�E4�A�~0L�|���	?����g4�Ͽi�N�Lh����ѷ�}lC�	F���q��'.G�]� �v�ͬ���@����Q�=Z���Z��;[�C#��T>���|6����E�f�-Q�����>4 Z���L�d���E�O�)�2�d���)1�Z[X�� �T��P��8w+�\x��Q�\q�'7s��R�WU5�r�RN�4�^�}')��~[&� �)	���~WW5}U=���:�5~F֚	L$}ˏq%�hR�-*b	�Ã}K���sK�Jn�G�ȑ!���½����8\Py�rH-���]�Z�G�fص_�qO��#�)��X�ψ�}sAV����3��Kgn��н���1�]1k���ˠj��e@޻��o&���]����� C~�Td (쩔��y�KW�T$�Uܺ��F��>����1V\�h�1z&Ĭ"�3`�[��	��r�5����;�Rܣ?�:e��*lC�g �o��o����������H�V�	�I�g\�YcN�G�j�v6�t5^��)��r�T�G�[�V,Bs�¨�Tn�(�H���BMZV4q���=�g��1_��Ńֽ��U:�'F��^NN�`� >�ӮABCsC^�F7BƓ�I�Gk��Y �pZ@��6rz	�N��䠆�=�ngD��UR�|p���lA(D/�癥�-��)H��> ����7�A��v�:_ê�$�}r��5��k�|��Pc�w)�jUҩ�,6��*l�f�t��EBӲ��,/�d=���v��I����$�i�a55��lBO��$��g�1��(X�a��7Z�c�- �5�	Θ\���Y2�M;��y�G�mLLÔ�����=@x18�7�x���������m@x��X��D�%^<���sv���3�� �+A}�%cA�j����ɰ.ӽc�+2�qXm���4Sc`n"}�u�R=�oσ�A1m�����t4�'9i8�]K�
H�y��)a�S'6A!I��,M=�t���9��v8ډ�����Q
���ְ���w���`.L�
����.��>kV���_�l���Hw\u7H�= �?��oQn�?>��'�"/4<1h˺M�'Q@�}��Hn;��)-���`�@F%us��|G�9�A�h�E40���ҳ�UB�,r�N�e"�W+�eh�lxTg~�s�{	�W
���<����,�00w}�򞻧���7�=z-��9n�GL�У�o��u��s^���3�!0l蔮:j�@g����eG,U��������s�� k,��H��%2ve7���`�e�����6�X^�@w�<�ɥ��)gX[�����]��;���x���_T#�W!�a7|݈r�u&`��A ǝ�w��=T��V	'�����
D����G:��4'���Eh^�]8v"t� S�6O��S׵^��_��S�h�W��H'0̣����[�8"1�~ĵ��B.�J��p���u��炬�:�S8�eݻ���ʋ�3��㪑7E��ZN�σ	e�T!?��[Q^��gF��]�\�r��T�-x�Ç�3�sR h�Ҧ�ie���6bp����f�d�����M,��@H{s>$3�|��c0���]���a<�໩�?���!օ������T��}�z�}�1�R��pW}+淒�'��_��M$$��|;�F$�W�-�}jb*�%Z�-�sV���%j
.U�hR~dz{d��"A����R�P�>t�~�񮷗h����KХ�1�ɴD3U4�=Oj�T�eӄ_�Nz�ޅC�ə�/���O,3<yYeh��c��^��3��AtD`K�D����O���=��X�w���{Z����.��b�&Е�;+]�)��w���1C�f�aFܺ-�L9�P��h��}���W\���¾�3��ka��XF��
�&z
߾6ӊ����˺n
�U�*�V��
J�Έ�#�[���?����"��ã�A~�F�m�f�d柳��}�'��a@�Vgw�5 u�vC�C�������W�fcnLlA�&{aш>o�j�lix�.b�;��ǯ��z\��,�w�^#L�t~=���F���c�Q��?�����&�w���T�,����%;C��"Wc��b�[p���T�
+g@�%~L��A5���YJ�l������
�q�Y�Un,�l��ʭ�����a�l�Ts�梍\V)�6��O��zD���\`Ͻv�_��Z0 �:]^�z�����U�s�%�jE6>�hO
�֙"0���ȿ&Ǧ�P;ѭ|�)�#�&��G@�5B<w|�
otS3�S�9e��������ן�}P���5i��,��3/x�gi�M��A�s�}Z�ˬ�\ۨ�0���s�/voE2��E���A0�l�+я���.˗���P�-��hIy	I�Z��Dh�X| ��xȲ>��G��*�#竼U�w���ɪ�#t.�+L1�$4�#șuhM(�[�g�>�,�s"
�"�];�?{,��ʒ�<�@1����Wg&މ��m��=L�G���O�^��s魇�(S��y����9�kc���[��� ������P`j
Z����^��_Hf���'�m�4��(Jˀck��b��V���&ξ��*�|\�8p������,���hy���E~ v���\D����J�����s,��&���#u�V[�"���q{�U�e|7��9�	m\C~�����,�Nf���&�ys�����<����.��ܦ��(��jY{�ov$6	�\'���:�ʜN6)0i�����YLp���$�f��]�tC��!���k��<�R9`�%z���tS�Nh����ae�>�J�B *b�p��3rF�^u��Qմ�]e0�E������Ӝ�hB�-9�@�8t�f�w�ӱl��.쉁�.��
�h����8B�r��s�+�o.�u$hqS�?���ʩ.���k�K������5ծjO���E�
�%`���� C�/c����9���^���,�XA=!���8�GR�1�t**֩�c�	:;��M���4�����?��8�U�jvw���b�M��v���<?��,�)�V��EE����b��>��=���艘�㛯KD�^�@Y1�A�W�4��;
C9���_�Cr����;R��Ҏ{��ˈB����Z��d�Dy�+�DW	je�#k{����4�F
?˯]/�}ޅ���|'�����4t��L�L(��E@���"��b�i�q%�/�aY���T42��[���#b����9Ԃ�ą��$F1e�x,�'J���zX5� Fn'�z ��b�$
@�Ol�O?Y�ܼ�Ԕq��?Ǩ5:�c�Z78I����� ~�m���r���T5��ۙ0�u�B�Zm�u�w�v��}�.b�|t �۞"V�MW�D{����;�ɋ�b%8�Y���:�2�轾%>��&m3�R�"з=VY�b����� Y��& *��ѻȴ
�<����yJnT#�D�?��P�dO��(ҵQ�[�F�͔d�^h����0d8�k��d�"�|��О^�v(f�v����~i��Ͱ�������P�؂I�8Ssc	�V{�ؗ�����W;D4T&G�yS��\�͘�*[�1b��-�ATʍ�� �,��o�I"�g���{���c[|�f��>{����J%��G����[H;y����n<�2	�f=U��D/��t��6��D>QfAxȑ5��X���p�G\d>��A�.sХM�89��_L{�>�~T�FVn̊΃u�fr�
 1
�p{@;e�}qj�I�(�!�\0�a�\l�9�=Jqy������H�_��r�H���^H�,�t,��H)��4���M�u�g`G�;��S�~h�R��F�B�ZoY|C:d�~᏿ݫ��vM�
�Պ�p��N�]�7�� +�j�i�N#SnM����G{�N|�1�%��p�p4n��8��&�f�p�%6�ވ>"k��bt���i�?����ZT�D,%rm�� ���Xj�VO�����Y�b�}�x�>�I��q�z~:^7�J�s��f} -�h ?KnCR]d�b�uӍ��Xɯ(��R�/N���i+�d&�ntp��-�S$�.�����~��L�N��{���E~,	>���8�UQ*�J���o2(^�2E&����^�Gs9�@m�J�.ӘLF3ZF=���"}\���I��n�>I֨�?ğjKR6G���V9�����hͶ���	k~��l��k��m��_�7�]�m���X�/�tw�5 ���^:.٢3���]�ֈW�5jBMq%����h=Դ���=�v��C��!�ׇ�j:
�	w	>�rة�
�[��i�]b;O��^KI��c�2b�Ҝ{�+EԏЦ${!%mq<p�W�˓�qm�5��$��ьm@��L�݊VX����W��P�j�m$f��aj���)��Y���������f�/+'�䮸.J�̷PH���)0<E{�y��Kuy60�Lq�*�0RźfKI��TD��O�6�:P���>���m��M��L�/��Z��ה��]+1W�yd`����5��|��x9��&x��������(Ӡ����������,�g��Р���*��P���;25X��ΐM~m	N$�c�I:��y�fv�O�<B�/�[�����,��l�������;1�񺕷Hn-ιǾ\wc�����9H�۔!��ww���1��!ʻJ�8���O~���Hi��� So|�E�d)N��r��/G��="��e ��7�q�`\Jl�Jx��b���%3ԯ9d��F�T��.�mex��(�ˑڦL&��$���B�\%$Qy^jn~��;A�l�ɴk���� r_[K�?��̆=q�ԟ^fm\�a���.g�l]�b�l/0se�o��{��+��=7��!B-M&��ռ<vP�������y��*��ߝ�bCzI��7a�;�����*OJ1;��_-�!�Eߏ{/xg���|R��)5�>Z��Ɨ�c�\_<ԃK2�d�w�.b�wھ[>�
�����܍�Z�v,a	���#��2#FCp9E�Of�^G��P���ު��}��6�+�_m���wS�g�1do���9��c�T� s4�=����o���nt0r�w,݁q֤��]_X�`�m4�;sգ�*T�$8ѳWT�ݛ}k���y0�v����|���p �o�~����FEi~=���܉����%��@�g%� L��e�t\K��@q}�uy��qjSo���'^w����{/:O/�*�J̅��g>�a����
V�/���z�bB�8>�>��}V�J��@�vU,4Ҥ������5q��]���@N����j�q4L�,�n2R���-�evoY<��M��y��J7g�N��1��ͅ;=�m9�=�5'G0��z��n�	�~�hh��ԃ�}3�����I�a�$j2ru�1b�Qr&����^�am���@34X���ͧ	���8$Z�<�K��9�K��f(���[ 
X�<{��+al���S\�-h��`<HW��_�������s|�v����4� ���� �"@�<C�^�k�X�_�����z�YQ�O�, ��|
Q�R�����%�D��wp݄L���/5|������_>��R��V����<W��oLT ��'�lF���M��xB�q��Co�[�r�m�ݓs����kyf��������z���g:z��=�!��\0�C^#�*[��Pu���1YÛ��RA��]{��i�W(�	�q��!��X��LI���a���~x�����&�"���`i]�PK6�˓�A��3��ܸQ������<.�h����蓶I�P�G1,���I?�5d<r�?@nU��0��r�a�,;|������^bW�v��B�tW�����fQA��2�����o�}nl��U",px�F�2	;=qpk>5o�ɯ]���؂��ʳR���Sg�ǵ�wxn��_��#�6=*��e��QǼ?"�'Iej���ߚI�K�:�z���,%����˽�؃�� }��-I��I�H�؞<����qw͞�q�>�2�1��h�p7�Aj*�G���: nJk��鎹
z=)B���l�M��U�Q	�p����d��#�y�QՅ��Ћ�8�f����V�f|yU5�̾�}���+���$��z)����7��ы�Qi�;료�y���Q-R��V�xq���8�U֑��\��`}&e�r�������ȃ@�m��>2����N�9��j�T���J$�ߺ��AM�0[iFn<^�W�Q��yW�������~'�.�/���(�F��ؒ�m��i7P{����|׏8���S���[��F"�先��b�kQ�8We���*�[��l�N�)c���&��P:��C`���.���A���Wq0&�A�PK����6)�b�]���{K��ncњ8s��\�E�
��D��mGԨ�I��|�=�D�4#��>2�I���8j���f��f
�0Hi�A��v�v�U걃��|��� {!M{;�n��]���X{����֞ց^�́~�H�v~kUa=c��P��^,�Yu�ZP�����0�$�Ч.|=�r�;��S(�U����$�u���R!����CQ֥��5]2�nT`��ė]�飆z�q��ϙܘ��"�J�V��K��ղ��}|lX��4�1�g���L<�)OZ�yuS�����k�!�����O�b�}]һ�:����mYEQ�Vqc���l��:��+a,���L�I�vL�ېΡ����GB%e
�'�3�e��|�*����'U�v����*��I���0.{��8ǜ��;��ZN9;�n|ƽa��@a n-�X�ύB3m��V����O?g���b���g�T "Tܲ�/����D~�߹I���=�=����s�gq�։���J�|����F�@Z9�zoqˇL'�B�����!!ԃ��_��u(�A�̘���q�GP�i���[0�.��*����܇�?��b[���Y7S6�1���h�'jcq�]^߃�;"��12��{TMΑ�"�fN��+b�(O�a��F�(u�5�2aX�O�zdKc~��j�̈��4<��EwY�qP'I"El��s�#̥}���;��*j�iQjgUب#@�̹��g�Aܦ���30�]� 1I��=d]��a�G������ ��Y��jS]��Ia���g����)�P��Fu[N���7�y��/���pN�����<}�����R17�(~�t�3��b�WWp���ћ"+�.B��nh�۳��Sfaa[�0�hz\�x+�q#0����?,�,����Z���D�Xn��/�Y�n	��$�n�D��~[�:��GF[������Kp���S��,�V4_�^E�ޛdmJ�f!�d��������F�hCA��½Z)ԃ��!�mv�m�;k��ۢ5���~D7���hd�`t�R�I�X�*uD�;��Z�$SG�Ⳳ]���&�z~@tn��4��IX�l�H��D�P�M6�f�p�8��,t�*�]����m?��zDC�?�N�n��]��3��݋P�Y��]
�H:�I�EaL>dM�����4�9�$*:[�T�-�e�3�+,��ubx��Z�}��� GǢ3�&s&*�]ז����S7y(��h�L�F�-����̈́��ۍ�%e&v!2=��[�q��c�*�+	8`�c�j�����ݷ�����WrB����!H��ܤa�y2+�iG��L�����ѳ{��'.�]�E��cyT���_�=o�7�t��G��5v�����}����f�h��8N�*�"�Bl)�.�v�=�K���J��b=d��1������T
c�ZW�K m�	�̕i?I�du�A������t"$/��O������Ő�v�(a��8�U<�g �*�{[��AU��I)�Y��\j���?��I´s���$Mw��K�uA���ڄ�d�}��s��+��Y��.·�~�&H��>�mf�"��M�]s�q4�:ߐ@�$V����W%����V�?tiH�����Z^�W�i��R	ũ0�w�09-�43��
�w���	�@<����h�W��sT(k��)V	���#��z����&,���E�5u1^:H��X �~s�Q�<�E|"�0�F�,Ҏ�{�BX�3
���f4�
�����u�;|BJ»)G��G�I��B�,9��P�\���
���o�S�(B�#�!��Ѡ.�?Wvђ�$ګ�������߅�j���ǘ�D� � �7u~�)ZDr ���M�����6j�qyLo�5w˾�sC��q����$��j��Y%c-�T'�X�B^���&ȱ3���g�j<N�_�9��Ib�^�l�<��!o��w���G��0��}g�>�ߥ:D�b�as=��A Zbh���zؒ���}y�R`���@?�򩭎܎�4oqcW�=^�5廘�_�: ���}�FXo�Z�'�Tn�yU����1��	�>n�G)�/կ�M�������O^��0Db=d2|��<%��Xmc�,��MY�r�I��9���M4��	����K�������	���}�!�)Yѣ��5v��CI���@l싩v���5(2�Q���5 �:��)��щnB��G�/{�0��<vO�a��`�U�90`8�$��(4�bv��ׄr�;_��mh��ѠSY0�N-�����E�/,�e�?M�@
͏�����?_��G�i��$���%)��-Ct���|��W�י[Ӫq��o$t����Q&ü�����o+�:'R���
���6����5dI#���6�$5֒c&L�0�����e��+'�i�b�q@f�m��{2���Ȏ
�eM4�FqNv*�-�4���og ��ŭ3�	h�p�CHZ65�ڗ�|�]���~���}DJ�����mɑTO�����ѓ�ɗ���e�c�k�*��k_KU��!�|�v��M��y��!��7K@�}Ʈ���-��n]SgU�K�H�5�j	$$�&��[�!(�g�>K杶�<DٜK@/V߁>+�B��mn�()���ݸ���3-V?��z�3@y�O���0�6[lȥ#u*�2Xh_�loԡQ�*���H,&?r���,��,��x�L�Wi���7Y�w�F2~�-��g�>��Эu�[��P@���[hWg�C���T�gg�IW{��I�N<g�
��ú��Y��Td�XƇ����{��?/�_3�odj�v�x�0Ny]#LH�4��
��咁s;��iݵ�_b/P�ݣ��H�|����*�����~��R@����0�풅>���(�D�f��`��5�}�ᵔ�>H��e;��!�#�5^-i��z�V��p��Ԥ�Чejf����=}�����gX_Q��)"#Y�s��X7�so���Nc��nڂ//�X�ڀȦ{��i]���5ǃ���z2�e�ȍ������1��_4�J!�����JX4ڦ��w"2PO��ĈTI 6kCm���9(����a�C!�E\3�%)�BEL�~���5f3��<e{���c����J�k� �����;f��� ��G� �}`���Y��q4\C'��m����i宯������8�4�"6A�N��!]̙9^[t1s���ZK(dؐ[����>��2�V�+��'��l@���h7F$��<��.=�ġJs�K<:����f[�cjd��Bx@��*2n4�Y8g������A5U��/��3���-��q�C�=4w�l>3����uc���Y�?��Imdq|S�M���`W�˅�t�����	Ց(���%9�E�K����-�c����$t�
�s;��Wb4�V���Q@k� �8�T"y�F:$��C��6��N�\��Y��jϬ�U��4�8����]�ϑa{κ	F%��:��#�3�\��!��T�&�:�J������J�[ h�{3�@�4�1|����r|WO49IȽ-'丵��H�텒@�R1zq^_�.��s�9S
�l���x8�}YP�EQʞG��}��k9�adϓ���1gBi.�x��<wO-"�5�Ӱ��c�y�d+,-�3�ޏя�q��3���@�� �Xt��MX�w�b��{e�V��j~��1m�<�Z��.��
�Q��u��X
��Y�.�zM'��b��&��L����7���M��\*�f:+�0�y��j����7�w8�I�eσ:�d�\���܌�g,�t�0����Ӥ���k_.�v�����k�ڣ�s��v�m1LJHL£([�������%Y�a���n��|�*���0�����z�q�d��U�,����ќ����{D��@ڨ�ߦ�$�� ��~��$l�@qn��)�z�T�ξ�ݑ����%����=l��!>O�s`�)��DFCw���9� iL�����P�x��%�Fc��%�T�]���NN�<�@�X��oZ�@#$��t �!n�z�[��o�*�!�N��r��#���K��,���!J'�C�����7%6�6��Ͽ�M쒨�)0G�����"�J;!��P�'���kմ�W}<]�Ɔ+b&@*��A�qߵ�!(�\?]Y�f�X�|�Ɉ����<����1�I^�l���Xת4��hK�����7��=i�x�A~����}Ͳ��&IH������C����Yp~΃
�������7���b��U��1�,�ި/T����&n�Ԉ>	n�p���\�sJg�i�!�q�g��ы�*��(}��d�YڳD�{!|jם��� mA0��.yY��)����#�:���t,p������w��f ��5�������vRd~ �IG�}���<�!/��fFv����#p�����\�ծg��W�{SU���-�߅l�Ж9h�2Ы�H���>S��b5�=8�:,^:�{�cH��"TރF���
Ș�l=�6�,�m>��N����7\M�Z����$P�z���:I������E0c<
�t��?>��(�$��~/,i��Y5\R�Nr1XS�3"�/o������G�c�O(��~���g��ctF���]�m[�|R�3�K��W���ŭy ���wFU��:�M��B�&�nFVh�?�N��1c�m�'�M��őDj6L"�=�^�,f尚Z�9Xމ�т]ޏE�{)�k��g3_2)�tX��!���}��U���k%yqWƧ��s˕�X��v�rNְ��W�t7�YZ{W�=�S�'���[��y�2��P\�&�5����bQn,�¯�D�ݬ��a��֩�v�G&�t��؝� �q0�e9ٓ^���s�[D��tB�������hn�=BB�犢c�|=�"\C��� [��؏v��>4�Xi7i��^/ӿ>zcHY�A����4$�`�}�]�Z�t�:3�X����vr����J ��$8��k������(���>�!�BF��[˨=I�7��Ön���ܡ� n���(�Η���r�k����V8!U�n�y����:�S��fP{b倴t��1	h�H��D����	�됝�$\b��M�
�J�Տ��v���{wD�@zʖY]b6B�D��4̻aea�( �U5⺟���� �ݐ3�8�a*�0-t���>��j�L�v��8�� x�u�i��䌅߾��~~j�pJ͟�1�`���0p3b@�1_��|���!g���^W�+*1:�&�X�"y7\�E�3*�lˀÁ�AUySŚ�^P�����eDfmd�+���	޽E}| �Xb�u˛��*�X�"��q6��l�Ntym+�sA�T�XG`c/�D:2$ΤñX�'BN��HX���'f��wL�	�*Hsn\R!=V��4��9�<�)I֤�}�re��U_�E�ܠ���$]4��!����p������=A5���)������2*к��p7,���)X�a�D�u�ƅ7X�8͇Hӝ����Q��#�8��i[e��\�܍OL��J�}h�2B���x���F�!=u_����a��.��V�K�a3@�c��=�[1P-�W�8�
��W���,���F/('Ri�����㞌�2C<ς��ض��t�I� �?�䱇
�1���5�Y��gB��z��}ћMg�\���^�]19-�`�����TGIM��i
��z��69�/%�f5T_��'���<]��v��!~�XLqTIA�En�8�/�~�-v�-p��\�͊:;?ns"�|��pZQ�q�܂�[ _�i�tHNmT2,H
jbD���������+��t�Ż���$�kt
��@'m��6or��.d���p�2[�C���J_e�ߛ������n��W�,f����͢�0�
��1�e��s��k�7,?z@�&)'l�X�,��VxA_�1�4k8�.l:��\���$�����+;�L�ڐ�k�Z�<�2;Zs���0��O�Z��i�1��F����V7�x-�0��`��~�o9!�w5��Z��ʕ�ߎ9b��Z�E�
�r���w?���ظ�iS���!e��v^>�w#��Y�mw��I�'��C��o�#A�jj��D�dS�W{��|���[�N����A�6���31A��H羚�8Lgz�{��C��������ה� W{�Eh��\XQ_�ac��w�z7�d0?0���}K�:6f���{�s-�	,8�!��Ġ��ӊ	�X�L��sznN(IJ��|y�'�+�Fu��#?{�kЃb�3�B�n�m�Ύ�\�� ?Xz��7ˑ�Z
��A'5�]b�I, �˹��	vF��Id)���Ҕ���pI�GmwM���`Ym+�J#�cf�8���30��|&�{p7g�z{�o������֯oNQs ��s�Yޖ�[GE�ާ�9(:_G�wA~�Wr��O��L֚F��H�j��B��� ʻޜ���S��Pj�_8��&u�.F��$g<�Δ�i����<�L���g�]��\
���I�'��@�uL�&�>��,ܘ����\�K��$�N!-� ��) $����W�-8�j���]�>\����s�%���b@��k&�dQ����ba��UN����b�F�N�.�Z%�:���v�x��'����m�$}�œJm�)�ZբӇ{�{�Y��������p5埋��Ӝ�Y; ��+��*zW2(>VSJ�'�\͢���0TGw���W\po��ӿ��K�Ud�]����+����W�s��<���Ae���j��	#�Rɞ�Rv��䱋G=>R���w�x�"�pmr~���%�����L��dO��^�㎂�����Q�GR��qּb� [��O;�Aǥyj�+½ǜDxɬ�j*#�6��T�U�o��@�D�7��0Z�����v�)B�	����m��g�Za�vUܛi�jL�k$���Cd4�'�اb�/0#�6�lmC��֍1�.yubh�f�ȸ��n-��+��ڭ��k���T�f��٥�:�س��C��D#D%%�'�u���H�{
L��y&yeG�.�5H8�IePQ��~��-0�g��Po��o��^%ލV��1QY�u�X��UA�H"��=.T��s����jV��'�'B&&�)�O�i_��r/�]��N,���Eio��@s��G'7��z�´zcN\$d�K�&�]��.��(Q���8�j�@3gVR�K�f���]uLT�W�j�R�F����@\�F(��q��7	�����X�|��'j3Ǐϯb��֪4��ύ,��*�	'>n
Qǈ*ht���J7Ek�j��Te�};��B,��9����h1D]&�4x�t�S��Ԍg^\�'*��-���d��E���~Iƿr�f�(�I��Xx5��TX�J� �?��ЧoT����z��?t�˾h\�q�~$N'rv�&>Գ�t� �)��>��pp�~�we0A�Ը����x��"D���H��ϼ��6���;7�e�="�K�(3b�k����N-�ii��Z�m��FŢVjȪ������P>h�z��ղ{��L$,/3|�y���0%īƇ�Z k	G����G�1�T���!�9p��<b�J�*?6��x�� #;F; �z�	a��p.���>a� ��~Ȝ\�9�]�Raex"���$��E�u�!��r�Xm {�`pj�M��ne�	��ӖC�@��"'Tk_�n�hS��u|�1O��V"�J�ޓ�i�����lS�W�ΦP�֒'����C�t�O��V�'o���v3���g�αppci �dwLҟNBޙ+`����;������EaU�5)N��΍����|y���K��^S�q�_]�t�:�:&�����m��iN�+����yJ��s��y�{��2-8<VVQ���F�(��iu2��f~/�n`��,�Z���:������-�\�����s��,���f>ov�UT�N4�svA-	����+_a���b�N�zd2�;&	t��`��a��$���������bw��>�!�=7�z���~X�F�Ф-��C��Y���A�m��4I]=�-�`a��Űzs-Bt�W��bV����,^�^��ʦ
��A�*�9ԯ��]nL5�n\
gH��?�����[B��@�<<I�d��Ŏ�s����w�C�)q �.�..M!1Q
�n�}l�ŧ��{E�Q��#�|L�h����Ș��ofs�z�[ΰ�"�Fbu>�)B�����_�hI��}z�t�Wv]8��&��K[��,�%�X'_���gп"�摌���o{3A_���F]�h>�ig�4F�2�#i[FJ�e�Y�AW����ot�cՒv��Y('��&��E#+Th��� �V6G�1���òj�o���g�m��?H׺DA��L���M���s!OI�H�&�q*.Q&m�1�O<�y���D��J����Srſ�y9�,��N�mFWR�>�؋U�H��*-ZE���HNosk�6�/n��v.�=L��Y�pL�i�V���Ð�u���>�8��
MtZD6QD�-aZ޼�C�N3�s�|ٍ�	�}A7O�����+�s�*�;��2��	�z���)I����Z��{Y�m��ob���"x�r>�.?�C��|m���1j�c��E�e{�7��OU����|N�au�owp�x.:۠����;��Zטh�P�ѽ�mv㸸[�df��I����.�
'�<ǁ�H�#O�#uD ��q��D%u�*�&��
\���]��L���"#@;Qa��m��b�-�Q����=x)RS��g���K�+�7������fN�l���@�7B�N<e��	����:�S���&K��Zg8��35w���/�Q=PBN�k�O�/�V	�;�ݪ����}�� �t��������(xQ]t�V�[S}�+�e,'ە�Tg!���*M	CT�c�ꦀ�n���^�"��ĭ8�!�$�rяA�ML1�-LhQE[�G��.��o��m���15���k�����1�=f�����e�d
A	5��Yi�son ���J��zPz5�O�m���ݲ����5����ھ�P�כw~vX��o�_�P��Ä�@�7P����Q��L�W�on~��fΜE�D���
�.,���T*�2{[�!��G���h�t^y���\�v8������uA��,^0N��B�+V$3����-� ��8}�
&YPTK��Ql��R�'ԈLD��V�&��HA<t� IX�2�=e�4�M0?�Md��CY���.�MT����h�I&x�lh�b% ��8���B�%./�n�R���v�g��xo̬�Y]t����u��2����.�	I��v�iHW��\�<��� �Ǣ��u��+�Φl|�z�r &/ �h���f�tҚ^��q��i3pW�߁�94����iS�8��N^S����'j߲@L�q�<�Lmm�L������O{,Ң����e����
h���W�8g��km(h�P}�^�^s��QS���i��5�<1KV�!�5���*'.L�!�,�4r�I�&Cxh�L����1Y壳���4��������宅��٠�^-�f������`?~q?0V+������Ba�T}�r5�d,�ՕV\"\io?][4X+��Hd|G�����[�}�rLb�i�;��qTu��T���������=�)yV[R/��4c����`U��*[�j������J��L�R/���p/����C�p.s}Ƅ�{�#G���e*�S7�5*��(��1�cW��y+�B�9��ɠ����ذ��k9(��.d��`O"��B�h������)| f�9;L�b��eIL�|�!`_`AkӐ��ͱ���'a��Q��V(��^p�Zg�7�m�� T�(�K��o����+��d�{�(�	�B�(Ǽ�o-�[~��TŜݼ�}!�hʷYz��y��)�v�����R������h���)$=wp]��}\v86D�>>;d���|�oZ�%��Z�� 塹Yj� �;����>���������4
�0�H.Y�'v^�:���N�' �Z���E�~������d��w@����T��7šj��K��!�]���K���~���{W�b�ʈ����H�Q�-0�`�0�u��,LQ��ԝ���k�
���`YI�����2�������]LT���1�5�&���!�C�@��V�)����8�x	ƻ�레��1 ���8��������A_J��N�|m�D �O]�������S�A��&�o�w�i�JNl��ƪ��E=�����%,��h�T٥�Isn��`�,
���M���Q�m�l�Y�����2����M�[mR��C�����F�ia]4SB��^�*��;��~l��3�۩,6y����<��լ��|j}�*�+y��zܟ=��l��H�h F�~�t�m��+�P� ]&t5��(��7`%~g�R�����o�|I_0��g��ęZ��'Ξ���'��+ -׸ގ�O���\�T�B�:�C)S(3�2q~�bB䭄,���I摅*����8�Vh����5����`�6����+��|�M�I�@4.��q;���%�� j(Qޭi����z�k�p4:����*5;fᅟ�����q�,�D�;�)l�����Ո^�b��->�:�]�[��$�f0�͏ی�����;���k�8A�2Q/�Uh��П��<�.�F��Eg�ൢ�Ÿ��#�(�łp�w�����YQJ5œBkf�wH�eѼ!��&M�ł԰J@r �츺�("B������yc���zF ��K�c*`��ӆ-�U��r���L���HV��j]�q�'{,o���C,�N�{H5��2a�p��$�]M�{%����<�@���Z6�y��ŕ&�$k9�������t&�����Vn޳U˒�>D����4�K�q�3���Ws8��D�xE��<��]�F�i��k-��<��5)CO���w�6�B��&��d8�cU{z�h���8[b�?`�q���bA����퐳��DL-P=�xW�0_>�g��8�p\ů�V���dgS��f������'���e�O{�&��4<Rl>Z+��[�i���lk�u'���ʔ�q�g�����D�����;�	��Z)Ak�wGcl'lL�iU��<{��̔TH���x�o�F�\'�V�I�L�z���:�Z
��v�xkQ�\�IV�B�e�J��BQR��(Gf�0��1�����6�*��]�,�+�*.b��?`ځW��+�ja�$_�fЮ�,�FkD4Ω���R$�~��8�����H�w��6>iʇ�=�HK��l��Q! ��]���+��IV5	��F�A��תm��sK��3��B�~I��޾&SѦ�~>�x��.����j�I8n�8(���V7@�E!07U�g�!��o쵍��c\�E�<�c�k����_����_ą#~�F�,f ɊH8n`�ĕ�{����2$�2�,���Uл��N��X��-��-�E���j��5���4���-��4��+��_;� q��ϿT�W4�����=�kZ���e�Pݫ���2�(���G@'9ŝĬS�R���I��b�gl:�"����N^7���d']�ڸ��G���hѯ{Y�}�"��ic�\���@�M�n���=�*��b���?p
��,�d$2*��RO��]�����{�s�a�|����JӃ|��=�SJXuS�/��9�=F\O�ng�uܚ
���Cb�<Qz������ ݿ�;!T�n�K��;MU� ��8�1B-���_Wy�د �U��Ɣ�)�_�����s�r��0�O�^��S'|H��z���'�n�<��~$��k�:@=H�;�����Glu�����������&��AI�}��K����6F��*Y[�Q���Ǜ��D�H�iC�,8\?����f��+{�t<�/e?��O"n<�����y1�M��"P�`u�^�Z:G�lM�L9�$r)V��au��]�	lK�\ʿ���?�r���m>�[�njo�M��d_HU���l�Ԭ�sb������S��[GR��N�X����Ʒ�)�ߤó����{�Y.�����J�[�b����.����z���N�=�^r[¤�t�&�u(WՉ�v�5��G�\儛G��˂0�T�ʲ	���5˿x�Y:�:��<Ẓ��Jү`6\PH
�#�vSc�w��z� N8�*B�@*q�e�|�*�E%k  0R��ǅr�1X�l�5�h%�5��p�M	-^��u�ߚx�j�o������A�E<;�S�Y�}�wn6ӳ�����0�5f/g�w1�+o��Zu-�s��g`�u18;Ÿ{|�r2u�K��-D�J��굸R���g�����KX��q6P@5{�A�`����Z_N3'�i�~�.�ǯ���I�����G���?����ŹL��A�t�*V�g�qr�k}��l]�BT&�$��M��v��	K�^�6@��*N��`S^�;�Nj����_�U��;����.��{�fN�PW}&wl��=�����.�hP��n�kP,�Xw�����T�
��x콙N���;w�}YW��S]��Nl�?S��������X�B������g��J��3l��x&6���A�OX��SUb�8�c��M�1q���������=���h��koK�mǎi%��/A��Y��D�_�ABq� ��%j�x�5V�.�C�����Ef�N�0��r�k��U$5�l.I_-���#k0Rn@�uY�Oyj1�_��<Tl���}>C��4Tz�)��n%�인��HS����#�K>Ck]A'�'Q�"��%BBm~	�ٺ�	yz�(BI���|�d����ǥ��	��A c#��b�P)�l�o{?�Ҝs!��ё�0���ṁl&#^ �
M(�?ǣ�q��r����<����C0�$�Qb�uw�j�e�~1�o@���c�^��B�O�ل��m5I�2k�0�
5��G�g�,�|PD�5J���h�5!�b���n�D������G?�t"�)��ȇ���_fe��*M��9ͽg8��QJ�<2������n�.��GQ	(�DT����PW��;�(�K�)�:2{Ϳ�5�,��j�jlZ�+�/,J픑Zr*`����f>�i����)�"l�x_/�#s��w"5�]��Kf�sh*~�ELL�센� �(�$�jQ��#�gdg����X/I�IL���8�@	�9�X����;������I[N��a�li['�Î �	�=��t��������	YZU<���mV�i��36�@���I��%
u���aS���t�Cr�O2��vJPv���q�v�^�o�}��Gb��S�(G9�w��A����)���6�_5�(-���!��+�;�8���d/�0�z�X���3�~)o/,v�~�|9��.����o�DÆ��Y())LC�j�	��,�t���FQ�������� �j9w�ȭ�;�L�'3�D���n���3���(��@Ɩ�D� �c���&Ҩ�6��� A�����̼���@~��ϝ;=?�P����x	֑������B�Vc	7:��aA�{E�Pb�����P��! c��o�Tl9��vn��d����3/�SF�<��O#f�6�B<t}Z"�|܄bp��7�r��J"2?4���n�98�uy���§;�g�^�V$��B
����H_~�P���V��|xU�i��z�3PV0!]�A�4DNr)"e��pU���ٽ�Q��7�7~��v�
.=e}����r��vHu���=/�D��n�[��
����b�m�Y��b>�#U��3BC�#QӞ'��BU���(�d������<My$�/���qN�̱'�Y�{}O��,Z�����$HU�M%�KE����tfPK6���"���5��V�E���9z���dР�+/}�y���ב���b�I��������SV�z��ǁ � �l	n8�)�O�i��wP38�X�#:7w���;):��\�d�D?R�q0�E���?[�3�	���U_+�C҄WNMxB�3�W�V���͐,=T��6���
��S����0�ۍ"T��l�Z���=�G����p�0�Q�~E�D��ܭ'! �Um��"&U���: ��i���,�-��HW�Ѭ\���a��.]'��v=MfQ��p�u�y��y�t�s}䣖�wA��.�C���3��5�F����7#0��c p��H���p�B��!0Ks�S�ƫ9��hM��\�����k�?��QMpf��q�_R�kl�a�ߍ�;���R}ӳ��51Wn����CO	���4����uJ�����a,.q8�Xa��1�ާZ� �R���	�)���X&�K�YS��7A6��I���t����	6+-��'�����_�	%�Lj��	R?U�<:�^)[
0�~�����t��c^>D9�'�r�1#�;48:T ��P�fXV�A��%�&�U���{s������%M��A]��my�>I�%{�*�l@���^lT�:k�AMq��O��B/z��K5����喵�9W	~0{���Om\�Us��P2�l�+ ]DL���n!鴩�@��Z���	�|,e�u�A���$g� ��^77s���J��H�U��K�Û�����`(�͂^+{���3Qރ)����7��s����؛�ü�����UR�S@3%�y�o5�9��xS�DQnɇ�7�l�4�7w*]G3o/��A��ݪp!��;*�'R��g!;<�-@���]	���N��3�"�KX)��=�r[��j�\�Q��z�C�Aw#M��hb����I�@XX��Io��0X�/��f�5�vPk���s0���K���g?�NOjY��[�c��?viɪ�O��(4y�O6F���zW%X
yj���~�g���q�6���h9�sGh���-Hp$�{
��>�?k��⁩u'ف��)@�-o/�g�.������c�ތ�5@��j�h������r�r.3f:n��ψ~���y���|��
�+�s_�w�ǿ�̄�M��_�����px�������y�^�:�BB-��C>��F���4�C�=��� uf��ﱖ����S��äkˢa���Q�Eh����[o�x��W�N4��}i�
kh�T�i�j�I*��3~Ǣ%�����6c g]��ލ�檵�7��Ct�oVcI�
�H(�|�J��;<���2�Wo�w�.��8�<��y�Qd��6�|­.5�X�9��,��p� `9�~%�-�6y	�b7Į&f#��@�!��̮��f�\贡1��&��H�~!�C��i-0$R�m�,^
�!J2��?�,��;V��@���&���_W��1�.�b�M���,|�(�FܽJC�>L�9�*x�e$��V5 +:p�c�O�n[1���f�KN�E���y�/�JNK!m�q��6J�_&v���xӺ�y��6�������ٗ�d�>�;�Iȶ����E쯝��*MR���`���6��	��Q*�}��s�M!�ӕ�i"��u��[�n��6��]�'������MQ3���/�(5��*��氟g��XPK�sN�O,��aka[�^�_����=V��@�n{�`�7K���.��g}�W��c�����5)��޿��.kʗ�,;����s[�8�D��K0d>��(���.6�_^����Z"	�2yN(�<�ȉ�3�R��j���+�-��6ɘYxp�g3j�a;X�6�$�II�R�f{7�vDR��{6<�,9 L�#�;O���*G8J�q&)��7j
�=�`��ͫ����8���ܧ�2���t�9Of��?�>��������?9�?�Q��z���ٙL�f��x[;̲4{o�R"�����2�5�dОD�����;�A��؉�8����Yj���&��H��>�)dZ�	s�o^�=k1�k~<�~*V�����n)���]��v�=!,����݂��ڡ������v*+T��_�Jhj!8�B:�>]��>EH�X��)ߚQ)�����(��YPkwGaݖ��p��!�ß)��LI��/	��_E:�/���w�35�y��E=���b�����6v�&�XؕTʯ`�0޼5%3
��	�C��x��^�,�kf�p:I#e	�@ǭt�ߺ/��#=�����x�'�b+�jSg%�d�4� C��aP��B-t%��C�i���B�;P98S{<������L�_Z;樊�Y��|����~~�$V�0�p�A�5��P5ي$��UuT9��LNI\i�SǇ��㕎�^�2��n�,�"S����+���]��\�gsU��7R�%�C8QdԄ���ݾ�p��(o�6J_#��ZZq\�ݺ�Z ���c�V�I��㎀�����0n���MC�4a��׋6�t���,2v��k���o��Cm��ZD)N�l)yƾ���n(F �Kf�8�5�Ks2��V&a�MNm�5����?���TVA���xa%���#�%������e�N9�|T��*EreCg"ކ�h_����t�e��4=)��w��ќ-7�2��RJJ~,^�0��-"�����/RS�'c�2b��B�Y��~����D����!�xE�~��YI�`�<Z��S��0����j,��/��w�] ��)Lg�o�Z��yY;T��D�E�@jW�EqH�O4d��ۅ��fr�*�7�ؤ�ј-�}��иop�� f���?jۍ_�!�X�tD������é+j�<@#/:�4�ZM�j�e�)�0�:����e�J7�r�=�O_��c�لX��NFûA/�ą�^!{��`uA(�S-r��	>`B����0R������`��"g"e�	�gG��`�1"�!������T��oQJ�7�K��Y��Z軪����Ř�EL˕$�@ݬ��Y��>��^*�j%��gnӽ;���ǣ�������x	��;�`� [et+��tp�G��A�L24�����k�z/P�g�C*J��D�-8��ԥқU��"��6fh4�sC�5��G�� ObVcW�-�L��]����B���ڌ����S���,C���tvJ���8��������T��l��G�^,`��֛_�q���!^4���P�|�N�(5i��?�v�����-l�)2���ɹ����R[LR�ƫI.��2IO1n���L'4�N潪��������:h�Uf����àp���2EpF��z;^*�D}�x���7Fp��:l���{q�bQ���zx�)u��JUJA2����
,�Zڜ2���Q�"D�
��#qa��������ӝ��y���	ֳ���Z*OS�y�{Ji7y;H������"Ok+d�b�#[�wvǷ	������,���`)T�|+��[�'�E�2����?�M������EM�������c��7v�Nht������0���8��!Dvn]��zC�tF[�-S�PA׹��j��m��fMb-;��ER�d�Q�f;�;E�,
��ck�6N��=e"~��*H�� ����yk���\��j`=��|����H�L���軏�H��帨�y����	-!�y�1��)��+S�#hw��)�s�ɢ����Q�����W�	`��i��@�a�w+Z��g�  ����fM�Qd�Z"K�<�7)��y���f����.B��L���v���JO�Z粇����ҥ�U$���m�瀊+
x��$�t�t�c}3���A~��rp�} *����l�=�_�s��م%F?��|���yJ{��w�8p��8>�C��	T�*�6jy�Dc�4���_G�m�8�7��O�h
e��d؞5?kᵱq��! �!d��l ��
��9��)����÷�5���%�+<���"��W����>a.��q`�X�7�>l�^;��uNK��8b��:@��ƵeuHI���&e���d��X�4��c%m��޿!u�`̩Ue���O
<Y�ysg���0���c�cJF���S�Ota�Sf�,����C��:�|���1�=�4k��7z@�i(��U;�����$�>���%6���TkK=���Å|4,hC�L,&�t:�.kKU�^��� kl��N�;)T1x�Ң����}��>��ߌ�@��сڟ|j��I�w��j
�ی:��, ���*��#��꘳�{2�/�3!��M{+��Z��P>�3�5Nk�TjW�S��#�}X>�X�Yl3S���!gړ�2��{)�����t������#ٲ��2�2t�/����8� $�M�&���ͮ#����PBaγ&�M[�9�UJv�7�}��ɔf����c��..�,���7�z^~�~�nU���2y�y<2��Ե��.�$��Ʈ�_�irۻ���?���{v�N��w�kڗ�:���@�53�;��?#��Ǡ��ÓT���~��\��\�������E�a(Z��2�H4�xbݿ�W���fji?-�����#`� �BI�; ��dUus�w�(��+��E��д�Fb0CL�m�M��12�(�ܸ0��s;���_.|$���7��VC�V��Af��n�]��.s��%W<� �I�ju[d��ӈ����Z�A�ȽR�W?tWF{1I�!-�̮��(x�`@�;D����U�rգ�L��t,��#aԺ�cbƸMEm<�:��BA���N�*�2�7��һ�s;�G����� �!��3K)�I����}���T1�?1`��6X�m+�p�����c%�iї:rC�/0�!Q�]�s���P���R.��G��1<Z��lj��FW�n��o�NMB���)sػc��A��{��iU_�.��A�C>!��E����x�E�l˽��B�d@`��;�
<�1Q7�0�y|[3~ȌK�c��tzp����o���'g��O�!���*����Z��uba3&�/�>�`�L�0����-E��2G8}	7l�!�@�&�+ôz��H��8��.1!��|;|�I�E/�2�;���6P�WԦ�]t�R+�L�]v!E�p�u��[��	���0�y����č�4����FLMd��w;�nxV^/���h�k@1����=T롘NAAs�:�����<��N��G��$����6;�ũ�j�Ef��Me�ZN����3�N��I�ڼ	\r�󃏝����� �Q�~pDz���Wi�jʎɉ_�v��m�(�$v�)A8�?e5�بW�����P]�>�H�AN�iz�8��P�X��˵�~���eZ>��ER�*Ɵb�>�_�_��ص�MS��	\ls�/�N�JʜA��B�!���ኧ�4_���X$��&� n�C$�vGEb�F�h�A��ђ�5p��@�� G����	6֌��q�����xI[=��[�v���=s�d��_�^S�v�Y�
�O��TZm��u���D�>;�N���<�}����QC1D����M��`8)u�c�:R��(��!}��/a(`f+"��˩�Aֲ�����.$Zרꄼ@1L��������E�3�K]\p���îpw
qT~}�V}�����c�[\E_	������.�����1yB@�f���St��o�l�o�� ��*G��R��oo�)M y�t3�7��n �_��� �X�4��랆�wC�����stV��0	z���
���X�<�:j�[��m�Z�d�",R���٫�A��a�q��ˌ ��Tr��R�n������%��݇��x���K�T	ٖ�ڧ�{�K��G��.������*B���R%�v�by�z�V�S�S	����Ņ��4��9�܅��+A�W���31�m[�E(l7���;����R h�R���\�CZd6�0R�4��S�Z�ϡ�=����ϟ#�`�ǈ�*�_���u���\�?�0wo.��-~I!��#�wC�F5�AĉstxN�ж'�v���Z��ʲՏ�Z���'��ʶK%`�E�C߾�������n�>�Q����D�
���l�����v(J�6��{���[U�g_��]O��3��Ā�B�ڰg�ܑ��X�Rʿ�jl����;.i�H�	�)����|gB����K�s:�%�Ke��B���~��o��:G��w��, �c�(���-hub΅#=�'�5Ʊ߳���z14�>�:BS$_Jc�[�@���H1z�k�� �b�
��L�~m{$����փ0	�3?��?4��7�9��R,��\��~h��A�ڒ��qN�ZLSہ��(�w�4��t�Tݯ��D��Ӄ��?�_�mMȗ_�h��:hC���A�D]0�!ܺ�0_�5h��'mH��kHvT���R�n&^�4Oy��r���r�]�T�-���Ѹ�X�&�;r9eZz��3$�c�.�.۾��=q�&b��/E��N��&�=�wQ��!��$��R澂�`�u�Ƞ�ITJhY���r�P`��	�}�F~�A�_���m�U׿=�/߆cm'��s����"<&���-Z��^	�ީM Gh�c#���1f�Ujp���͔�u����#L��Fy3��(�+ȟ;稱��w�_�"�xG� -�ͽ�V/
���T0��+�Z���K��H�mu�	~bCBY+^Ӡ���eSGhV�6�&dh�]ǅ�z������Ҁ�<b���;��*<��>"��D�.K�\>R�z]�W�Vsk��`7g�.����>�HCFv��?�'Z���>T�����s�&k��b��.�� ��̎�m���ZV�w�E!m����,:b\\n��C_��
� ��ǭ9�_���O1B.���4rRL�bO�c��ݱ�|B�AR�|��(��D��� �]EE#}��5�AI)�U�B�l+Y0���-���k�j����E-({ۭYQ��[Iap�^��Q[Z\z��=��6�n��ң��Q���Αn�@9a̣ C�7?f�M�Qn��]i�t�O�x���T�۞z��~g�6�f�>X�ܣU�Ki�yѶ�m����d5&J+��8?����͇<\ys}��a4w'�w�p���CmC�{��(��bn���0�%��y��	4Ҧf�2w�?B�cy����5��TaǞ�$��ɹ􊸏H�C�h�m �|�h��*;�O�tpE�y�f#���FQ-f��������������+l��-���m�yH��k�<�7�~��R�[p5��Y��c��K�?\���)+����ɦ!+_���s8		�����>�0Y)����#�����_���,��k�_���2�'�c[\�5�e r�d����:Μ��1颍2r�An���OZ�.D�w���6֏й�7&���}8O�W����rL�BC"�]�Ϝ�j:,R(N�P�Wِ���]��*Fe�������1S~�'#{yU+���6G��!}hv�gʨ�C��[�V���8wآ:�l�r���|.��D� �3����U���T�5sQI�U���'�^n��%��p.!��o�O�P�s�O9���n�+Cn����X�*���'�0�hr�b~��U�Ѱ�r��ܶ���x<QS��Ҍ�=��H����`�!%���
��y(cL�"I�����)r��QF}��Q��>��sQJB���;��7�Xnj��_��jU��	7-��l�g�xM�b���II�ɣCk�b!=��R�]�0��w�ab��j��g�'�.�$�����o�׳��ևrŌ٩aW�� �M8���o�m�8ꕓ���=�O�F6N})e��U�	f�������(d�(�98��a�|CO��$�.h=��2d^8W0+پ���8�K�����,���A꨹UZ_�D@�u��b��������C��W���){qA1��~���T�a+�������GV
�A�~� ������Y~��ؤ@�g�
�ը��l�X&5��'Dfx		s�?�J�v��y����TnR�h�{�B�YZ�k�g,Zx=�'���ΤiF�0��p�d�+�g�a_�gjb[��e�4]^sqSJaG��(H�|qV�f!C�`�H+�w������+�.0�l�vni���ȶ��'�4��H��Z�����Η��K�+`��ɵ�B��B[X����2B	����wXW^��Z���-R� ��idK��N~�Or-VFs
7��IM�G��{^�'6ʽ�RC>T��A3~�t"��_������Fٕ�u� ����(��J������#�O�G�D�TO(��Qą��bjk����vCRG b�<�
*����?�@��Ռ��%�j*��s9��KH��4l��9/�g��i|�Z��5�-H���Q m�eY�M���sg��ϸ�I��8��]-ID���|����R��ο7�gćQ�]��}��>5OqC0���r�1⹙*>�����D�vk!u�Ĥ�.Oʜg�%��}O]]}�o��9d�XV������-HMk��חǇs��E�_K�_�Z�7g�$�ji�� /��j}1�H*$�x{D������	^^.~]E���x��J��@��؉/H7)�,�9��n�׫�-$'?=����q�%N�8��yq����� NI������MA/ �}�M\���H�&����4���F�\�q҃ݛ�ߤ�hho�f�1־����<��o���P��$6�Ϸ��M��/i�`�*�PEv�(�k�H��m�Wv�h�/�A���	߲~���:���Ǻ���g$C�<I��$�#��`��rl�#a�kGC]J��<Y�rB"� u-��z�J[
��9�D�e�Jx�5����}Zr��sz<��1�)�)�x[��R��hl"`�/+!C[7r���*�y�F��a���.���<�L����X6a���F�Rp�z� 1��fw`���Q`
��0�S?�<Y+��q䈠�!i�A{��{V�1�݇�@����3Gn_�"��ֺ�z�Ù��Z<�Ӻ�Z�OPV��������ˀ���h��8:Z�܊*�+d�-�t�x:���|���v�� �{/6�᰹t��ڰm���E�N�D`�"�M��Q֟/Bs���� +�^��C�z�:�ꛋ��������GB^86O�-���)D�}��t&�*�Q�/(iA^I���ٝFX�`�� �	�ɮ$���-b�d��`�u�Wa^<�n8ښЫy�G��9�ͼ�QP~�b�5 oEP�6Я^�Q���q���+�3���t�W�ص�\0ˑv���O+�A�ЬR~\�mő"�mU���.��|��2T�aUx��k���E��ЧC.9G�&�P��q~p�y97ģZ_K�,�-!��a_ �Fa����?D�[�F��J|{�T��l2�JlF�����t�:��ʹ#q��{L,;��Mm�Q��x���tV��8z�"bM�"l�&t�к��I;@�����Ǩ���8G�v^_uשOƾ�@��D�ǽ����>�d�q'p��Z@TI�$p��d~�E�<��s�'�SOM���7X� � �a�2Ƶ�#������J3���Crt��O|�UYe.��wk%d[2��0�Bo�ZQ>|��k���s�!����.�'
�τd�ݿMG����w����6�p4b*�K��Ml۹_h)SGc��mⅈ�p��B�z���g�9�f�BZ��GV#�JT�ט�&��)�����'����$D��I�C[V��r�|bXl��C��0��]
x�	�h�K`ҫD1�
Q(N0�a��D��I��AP����6���Y�=bۙu!�3���W�L,��G��4ͩhb} C}�Hws�1���ʲ��ڤl�HD��D��]7�p8�I�?:�2���^��,p�I͐�u�?�x�`_M�͂�a�>���ʽa��"��~qY��زȈu=j����_�ѹ�uF�e8�(gtY-�-1�����~�9�F��AU���;�)h�eqs��9]~���c�ʾo�3�9aS��<?���Ɋ��^M�+�q�SNeY�WS\?O	�o(�͢.f��UJU9�=W����׃%�GVTWF%��D_9�eZY�M�G�S`����	rч[���e���&1p�Wa��?˧�O'�<8�(�֕���b����O���"N��(�h'���&�(0����K�������}�',�U/ũe^l=6��_�6S�ܶs@�	2���"�h�Ni8P*J���K�
5!���umC<��T���R�� QK��*����о��Nj���=����D�_���a$3p� X�R��_۝ N�~��@�*�c��հ�i��,NnC2٠,���cٸ�}P��W�wM��Ү���w;��ΎD��?�̍�+l����t��e~ ��Y�x�����I�(T�z>��Hq�9�M�6*�+�����1W�hPLi�y@�w�p�?!�o��^�Gi���'j$�ׂ�@RoFg��"Nx�|i�0���êK��F��~�1�{}�זø�l��_3wʪۯ^"
�_�W�-y]p>ƫ��O	����S0>Z<p���c�ύg���z@s�8��Y�-�O��/âƉ=L�M�au�Uk��m�e�~`�ɢ��1|".��jp~k�X��؜�	rA�w4���Y=_C�U�/�W�{��������j����Na�}�u{��1.h]@+���h�?��紁�pO�eM�	��`��T)	�w:�2-~Y����c|˼��!�6����F!�N牆ǩ����=�딢�־[�"~�ŻHK2������b�f0'ƪbn.��.G���4`b�w���6�6.U|��j��]�j��<�v���'K�UJ���M���ؚ��r�M���"�fϙ+*���;�[��l�e]�V�u��o���}^��^��� �������I�՜8����ۘ��&~$�>���C;X���a���^3����~*�`I#|�#�|(guw�`��&6��s�/J���ͫ�(`���� OVmy����{�
$i�N(�}R������4��.W^'[���3�V�)e���u�o��Z��]�?�=rԔ�Y�����~�0bp�M��`�rx*&_���F�ю1{�R�HC��ӏ!��;��z�Xo�k����D����JX⚋Og.���۪h�d7��bb��O$��_�!�q�9r�+�%��� �_2��~Y�iK������9�ƻ>ɍ�@Ÿ���׀ѱ>-����=P6^�����n:�sF_�iB���I���� d�,�4\�z��+nE�����D�ѵ���㳫E� g�N�7pOi�O�� k�)wm���<-���A$�{j���6��!�~�f�XMxgI�i��B�<���]���Ֆ�Ǳf�ĉ��0�g�xh:}}F��V��l��T+Jض�Z�?z�>�v���2�����B���*�U|�N<�~�@*�[��CǷ��1��%c"�L��U�u+F�`�r����KH���`�:(��)|�Aڹ��3(��!�;RQ�qV���ܒ�'�6�3������SX�A6����,P)�U��sϵu�L��eL���V��B&���x�&(����
��`��и,����14 �1��z�����%(�-�*���	�;1��p�}x��������:��cWt�q�j懒��B<<�P�|/؜�9I��Վ��q��Ί�Y��I���61�:Z���*�OZ�]Hp����Hݩ�'F��壴1�O�]��A �����i[F��vl�Z���,-�%i�NVk4�Gh�����U�#-U����e����d��̋q}�E�k�;~Wӣ�D�V��9J����ǏO�F��気���_�ү�������yȇp���d�M �Z��\�K�t�B��Y9V_AO�J�{B��M�ȻO�6Sqo��g*C�'x{�9�RAPHc<��\����hf�V�����]u����#P��©;�P�ƞ]z����^��V+�>%?h�p��:�����s��-iv��cFvQ"�0m��X���̑d�\���G�M�~�{�ߖ�R31�S!M].0+D�f��x�8��b���߀'wi&�0�w�,+G�3��{��DVT�2�O���-w��z?�7��L��2	Dq�J�i>^Љ�[����;���e7��:;�*%��t��[��-Km��#ؾ�Mc���cɑ��ŷV�?�'!�O��='mV5a�i�+��=S�w�Y���� �y0�5��on=y9��wD�]��('gϛ7˷�%S3E�S��#�]����3AS+9�]��%]���N�Eu>#��k�������DWo�����1���oR���~�3(���ƅ`]^30���o���Y߂�0y�z]��~�|#�<��i:�<Q���'�Ž/n+���+A��" �A���u�9ۅ��ۡz{ �:���b:�bV�/mv��d��y�ܹ��w���>��W�0,k���EEO�D�c�NY��x�s�Ꝫ��V8��"8��#��,]�^͚�{ň��Oe�����\sT���v̌�<�����~z�^%H�pm���PO����^�R�g?HdKYz�~9Q�Q+-����uMh���֫,7^��V
\�����a߈�\g�.��B�hr��񯃏��&��� +�O��:3(L�Y8Xr(��4f�"���+k�~�
z�"���A�$Ҕ�yBE-j��c�j�g5C�#Ȝ�f��dk6U�ɤs��_��l��9�(��_rI�G.�l�z㹩��yBk�)?��"իN��
�~!����i�U�ń���!���������EX�D��^��t&� D7~�Ŏۢ,�-`}?}���]0���OQR \�
QLL����Z�gjJ��)"wp�%R-�9���5��
Tv�=l���Bp)��`�����-i<J��r�:E*�M��R��2�$d>o�,��w�QAR�:(j��7t�'h�
	���r�"4-J�C@�:����2��k�ղ`2�����REY�Τٱ$,Z�@,+��m7�tT�K�ٻ/T�8Sc�������7�9ʏ*����K��O<C����S��u���Ǩ]_4Am�u����F�n���Qh���Q����x7��Z��4�o4�{M���GF2����W�5����d�&���\P��$20�v��}fϰ�ߌN�4*�W�2^�/�@���\�ޚz�B��R;�,0�'�ZQ��5���I�C���C�ь��`��6���c��J��*P�V��C�A4�^N��oE'�s��L�;�dk�zT�Dv��6�k�4"˺�[��́<i�BY�J�L?��I��)J���\k�^�z!���� 4��iEQ��&�Yޱ �CcFFG��U٢K�yi|� �L�؉ON/���Z眭۝��p����|ȡ8w�(�xD��2�	�T��?/2��� l���FX�~Z9�;�[�E$>�}�e��^�G���{���H��>1��S詷�����:�-��3�?���p����s(݁G+��0C�"ڹ�����U�䟪�A�"�QUO����?ƼC#���Z�$����e$Q�F�eX���Z���nIz�"��l8����0��_�2�'1ڹ��,�Z��>x-�0 ��(�)J��7�`4L�qL)S�ǕUD�<Q�} Ȭ�M8�G���]͑<*��k�k���Л�W�C8ԡ���ZA��~U����� ��5�9���� x��6���>�f�N��Ѕ098B4j:h//)}Y�b��lT�� �U��ڥDVП05+��� �ڌ�\a�-c�	^�Fvo��W��$,[ӬB�!歪���n�L;�Ts��Ze�������S�9B��i�d1����Dg���d�/��ד�~�b�''ΦrI3uR<�+M�u]�N����+rјI�����e'ϴ�	>~�[Z��!�|��Wd�K���G�&>�K$Zy��Ν�(�
`~��f�x��r�ڂ��#;��~�7�41)1;-��$��a'��u��q�s;�ǊZX�/-vۛ�k�������h���*q���G�% sx�%�qBߨ�a��Eh�91!_���̾/��Ko�pQ��*B�������m�z3�q�]�a���|;�L���2u�L�)+�C��yd�j�dH/�i���Aj$�d��q��[�"��!��� f��h�o>Ɉ�FX�x0)����c�H�\����7���i[Lc�~��|t�����p����بZ5�_�V�F0�;�%��[����"Sm������hYp;Rպe�jb�qO��O�w]l���T(I)2�?��{LK�m��
���{��%�;;�dBѧ��m���Ć�I��q��*0G@[=��X��1�%y��E��r�լ � {X[��i)\x�ml-_�f�(�R�����}Ln!׵)Z̨lE�yWi�{����׸���;֟.^��2���o�u�t���ű�l�|���W����!�����ѕ��^�ߣr7���)�7��~y��7Z���ك>B�.cF���)ۋ�4ߌ;\�D��%M�LJ'3A\Nï�yDKb*<��hojtЎ��E����!'^�`h|#��zД�J@���&�TT<p����L�C���I{Q�ZQ�Iγ�t̘Cr����Mߑ�wr�uH�m��ɑ�=~^���}~��C4U�U,_�Y�,��Md����9�邤�20-��̉Y��v+x�8
B�9~tkW懝O�N�4�����+����ڕ.���č���G�A��:j�Wo��ٝZ���&��Q����"V��?�l���*QZ�R��t�dp.�YQ7�V�6:�)v$�V9x���H�k��� �W������2����Eh|��xV9jR[��A���ݲ%U~�k#�EV����b0Cù2f<|i?'�-�� �F����F��:���\��G6(χ�����:{u���mQb��fkyƖh�P�C�O7�#k<O+ip��R�|t�a}��N��
��c��쬪Qeju$}��D����p;q�����'Z�Aʏ�=��mzb�oഃ�f��CX�$\Ǝ?�ά*\�������K���Oɓ�XƊ)�	!����Fn(�"���A��L}��18]W��8\�������й�����3�~G
���f�������{&6*�)u�:��9���r<�Rcg֥��9�u޺i�ů���$��
��؟�r'�����ӫ��h.�C����ɜ��_f�Gz\�8�z?\Ԗ����Zf�(t�����=h��i�~P���df^0�����(sY�M�*�r6	3�e��):+��a3����>�d���|��9>7�·�4���8u�7�F�G�/�z��̹�핃�� ��枚E>.� ^�����}�|i�g�]U{�B�,h���}0_�oW3 Hj�:I yH��7�w�0���|C���$��!�m�
��PU&�\��f��MJ�lc��p�p�5�C?
LqQ7|w@�T�"��P;�O_۔�9��nF� K,�VzF))�r�@.���B<��!��7vP(�ğ�4��<�v!^��r�pd����#���c�#��W&��u�A�Z���7[��g��Sg_CS����y���#>|zf|��N�8�T9c�@%F�>��S5�Y?I���Y�M�����]TA���i�@��u۸�d_X����{-rz���1 [��L%�U��n@d��1�& ϓpG7���]��-��j��p�
��B�T`�8�cnH�T:wn�w�����/�jJS����k�}j�x7�͙E�p�$</���$	�Π���
�3>3��[")ǋ.���IU�*�� 7�����K�e�`)�
�c�84�)���_�=	�p.)E���a09f
a���Ʌ�����JTA��G��2m0L���f���B�Y+�,�"�3���}�P ���W2("�$�5�Ky}X�#!�uPl���ϵ����	.~ۚBqV�Z�8c�l�n!$9����-� �(ҡ�a�S�\{h��m����-�P���k-'�O��4Ϲhf�Ų��Ty�s�L�a��,o�q�Z{n��^�C�>�I�_nq&%-X!vF��7�>L��Y�lz�>G=�٨�R��H ��Ϊ���E{^������8������
ҜlP2H����'�Y:��r;���f�O�aJ�C1�;^���*C��(t���"�D�/0�������Z��i^�p��x�Zv`���[����!�2\�ɘ�eIRԡ'ܨ͚e:�jW�f2c;����Ld�=��&PJJ� ^V��d�,��Y��\u4�edn��	�C�{5<II5�vj�[$�$g'��b���]R��s���b:9��x�_,�	8�lN����Pl�V1�%��j�&+×!�W��9���0��-�n��l}J�GN���Y��4��FE6Y��2�ak>�"k���yn5�0� �Ʌ��0�bg�� 0��Q�,�����'��s6�WICrT���{SBS����7�G��؏�_@���� �y��a#��S˃6�Ĭ|�e^�`���~��o �r�s�Y/����C~�O��H�l�Vګ�7���+T)�U)f��7�y ~���>����gv\�����p�윂�z�E2�6|!7m}\{�(i�w��ZuRg�q�����K��s�bug��l�$��d����l��kS�I<F�� � ���9iV�N~t�d9�I����E�j�a���uw�3�o�J/o'P���3��E�K�~�{:E4���^�:T���7�n�*/����qa�ɛ~C]"�򑪶6a���a6�/�0�+M��q�����
�_;M�S*G��J[�]�H�Ǧ�P�~���j��*2%�2Py;ª���w�@SRd�_	���ʥS�~L��d�I�79Kxֱ��∐��|&U�㷝���M��qv��7M��|�v�5����Qf獝�z.m�b¤�ovЕ"(ߌQ��葩`�X;�V2Ёq*��w&>�2I���C�gD����9O
�@c�Hp.�)E$��<@����
%Z�,�v�,kG����7�yF�Z0��p��\q|/���gE��^~��بPx�����.���X�����J��b��R��
#1l@|6η<5�� UTj�D�7iND-�r$��[��h�^��p(��}�,��I��o�켗e��Bd΁__��&���A�
��$����5�2�	E���������yj�JË��ۧJ�(�'��T#�h�Ǵ�ݶ�$W�ĔD�n���t�з�'���;��>���Z���j�쫆�yt�'Inϓ���$g"�}�r1��d3�j�Q^�(�HR�/��M���\�1vއNroL�h\j0��#u�p��\�.��H1��6��V���dbm�����9Yg���R2ǗK\�s����|��o�t����=�G
'W[:_rQ�E�+-;	��G>�,�l�Q���@d����D���`��@Ǜo/�	{��X��b8(���_�8��ny��������6������*�^���,*����Fuy�Jˠ?����;�ϑ�'�_uk��5<cUnn�e��Q��4�K�6L�������4c�IzD�W�����LAڍFx�d߱��¯�~�l�A��-F�M��k��]�Nf�*�4+� ���I�)���W��r�ǿ�ω�qk��l���w���e�������WϿe�4. Z
�^D�N����J�L|������k�0�k�v��%���C�F�DL�z����%����ݲ���O5)�K���"i��2Q��!��hW4&?�f���+pt1>�h�u�Z���w�Sp�3I����A��E
��ߩÊ�X�݋�7���qv�0���� �{�Ũ�4���0��g�AazU�z�7���8�'y���S􈎫u��>��]o7x"�jZ��Y&F�}��fu�����xrъp8@GMZ�e�~PQ�Z�� 39r�Ks���09��:��� �}zsGD�O�f[��@gg�������-V���$��L��f�|f�7�!�	j)��*OB�a�#����Dd�
�]S�M�V��J���X����N��}�~�)Xx��I��>`s�l��R�œp�p�7*�`ٺ�"q���|���ғ�� ��K�ܣE8L#Z��BN��;V��T��P�І�1]�^ihh�Ŵ����5�,�i�d����ɓ�ǵ�c�gi���'�ohj���j ��z��c��Y��P�p%!a�m
�M\�K�Ð��z'�Hv�R��L1c���q��p�:���,�* �5�P4��|��wa2u��/۩��F�	��Ch&xj��� RY�t;�*�q[�9X�4�.כHY�S�O�"�˟��E�#0�nX��ޅ-�A�I(
���$�ע�nF5e�8~ܓ�u�FV��A��Ʊ_�Wԋ_]Z��.����f1�����q�h�Nr��S)�����QUJ����>��H>�4��7�î^�B��|<0��Q��D%��^��Y굕pԔ���k	r�/���վ p:��b/7JMoUs�����E���q� i	�v�:Y���XR��D`�����sB��ѷ�!��Z^W����d�_qs!R^��ʷ��	�a/�j(���Ҵ[Nɨ�46�L��JƄ�S�[��j3����6h�?s\B�������<&y�I\��鑶��X�7V�F?�"s��R�i��c��B��%�N������e�E����GF�ҧ��X�v��ާ�m�-�1�sZ�*+��6�7X��c���D�������w]���_K��u�<\�~Y�M�!���y� c�{Bz��q�9��k|;��T�ϒӃ�MYt)�FO&^�����0�q��V�{��[D����%��l���V&W�A~H�k���kSDx��U��a��恷����BE�W�Ya�_�#o�+vTH�@=�WE��~�ݽ`Q3�f�sz�}����+�/��_o߾*����Nh6:=)n�?1e��O�8�~���^H�c�B�b��n� S�~��v�ndg��NoSs6����s<�,E�l���H��&|�kL6D�T�_��B�� .��>��<��|) .N�>�ǉ��#a��!c9���/�����m�XY�_4�F�f)�H�PRl��AV�b�^X¢fv:��sB	�C�b��u����M1�O�$s�����Jq�(g΃6{�N-�em��ed�5m���Q��j,����c�ټ�i�g�G�r���`57�hč'	� 砌2o���>����N6�C�-���!�UEP{���e�`�U#ul0c0Y����A�- <Z�!�"�o�dL�^��:���>���D�$�Hjs�}I�4O�Ύ��KO�����g1��AM�<��+��[�QBL�
`�\x&�^�Fd<5z����R�Å�|����4No#9���K��Xf���5�Ba��jN!��O�P����(�@���A���5�U����V���q!�B\�5�!K.����J3B���'�n'x��%zA�������,!
���M�L��o�b��5�W,�a�v�rf>d{w4� pa�a]ƪbGwBG�Z��͚�h'�FX��^�Y���v/m2"�s�p3���
�W������e&����!B�nHw`ꃛpO�+��jp ��kń&Zq�"0��o͇iP?�ɡ ��t60�����
P�:* ��%�����[�ߘ�1c���h��Ow1~F��Ce��_�AH&H�)�`�z{�
L���&>I�.h(�5���e��KKu��-rUie˙���~�"��=U���8$�7a3���̗��YpiUuT��6���Ay���?vX\&�]���n�^Sz���D��dxs����?ovq%%il&uf�wj�wz }\>��td��݃$ =��i!o�vX8�_�S�Y���*v�;�kc��E���SJ
���Ě��S#]d�k?3`m+
ZvByb�П⡠N|�'}ѽ��=���f����n�-l8��ȧw!tOP	��M
�hQ�
��#�Ӟ�b��H鮲6!�B�]i6':�X�l�m΍��l�qRg�7���2�����X탧�H�����d_xjH��FT�zr
�vRaH����/W��2��}Jf�e?�#*�� �ɿ�z�aH��K9��+xh'/�.	�3�)����F��F�V�j��$����L����Aˡ��p�&�� �d�<��-�2��B�t=UX/�\3�
�Q�u%7���٬�EY�!�&� _�X�DC�i-�W�6pZ�m�*n[�k1Ҽ���%����z�"p��	��\�����})w��X�c��X�b��&���1�&%���Z)��Y��p�!Ƅ���	�ւ/��+��Л���i�-y-��^����%�i@:0����WVg�$���YZ1��m�A��&D�:�M�|=�.�I���u�#ԨX_l{#�{e�sT�)�2W$��AP��D?M��1�;7t(�"�H�3Ѷ���������ڼm�Dw��J<T���F�"����o�r�as5����+����>*�PVz��B��Yگ�r7�2�i�k�җ('�AQ�Q��Lb���R����j���]A�!A��np۴����5����eB�
�r�،֥��ȗ�b��S� �f��
�-����Ǘ�u���
