��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0R��>q���Q�I��	�B�R�"w8,�zpD�ߨ�Zѵ_��jq�� r݊�+UuIǇ"�c*3[ ��BO�D��ǭ9���Q�:5�Mcrq�V��Zb)��;��{�|��C�u���_��ɒ�&�	:b<u��piw� M�=�?�aZ��q���+A�5~r��� �A/��&?�����W�����z�¾j:��f�
F�D�K�E`�j�Ai��B���&�WE�t��?���u���}�"	�����B4��Y���ϴ���}Ԙ�%mlҦ��; P����anE�5��f� �R&3��s�3�9$�h���/���k�Zq�E�U)�FXK�皾}A���R�pHӡkq:}�	=��i��:���\�u��	VG����_:�5��z�t�4l_�a\z��J%�7W[X�@�	�8�$^�P��-�s�g[ENHK��o�f��-���j��'��	���]��'�_��h��N],��������%�߯�;�ԴЙ)PUq�O�Tn�f!5����5c�Sq�=Ţ�!]]J��̄}�&X��(*�(\ |�|N��Boτs���f������y��[q���(���O�NJdU��^5�YDO�8}t"|h���q��8D͒��I/GD k��=jد9d�� Vw�n��˓��偘�ψ�q���)(��Cb:���w*�m/��%�b(t{��^�ӯP�M>��^�	�}�]��n�j�.?@N;��:"���n�%��I�fF�9�2;�d�!\�{t4I{��c��>��U�Yթ#��(4��Ow3K �ָ:�vN�APe��pc��}wq?@�orF��6����ys(��=�v�l��=�xs�c[/�gD3{�z�j�p�x��{[���?rs^�aa�[G/S�����T6�84�ؖ~�-#��B��g��nܘX�VC��8�b����?O�P�t<�
#`A��;��
�܆���2'��IK_��v��+���o�mdl���D2����؃��� S�(����ơ���b�T�z��>߆��]��45D;��������{���v�0��yH�U
~u��pAA�o�|���DW�Z�Ӆ��+�3Y���]���탸�Me��*v#r�)�ׅ7��S�m�a������4�p�'����G����I q�?x��C�%咱+:�Gj�˙��G0g���fpQ5͊����+]z'���d_Á�ۘ�ҫ�I���B��##(��2�(R�^DX8�>W�����Q�U�Seaֵ0MO�]�ސ��B�򮱙"��@׏ȩ�;a"y%}�\��w�%��62x'�`��$.Im�^��8��;�c<�^�D��O����mc�KV�1e��,���[�#�ɻM��.�7~�s�o1��M�������1�	B���!AB2__8�bdJ� �ZA`�/8� ;�,O��J�a�ڏ�� <��p�*{<uZ�����N˄��C�ӓ:�].G�m��8{���$%8)��������J�����@��C�@���{�2b�[ry�[ ZxP�c�h��*���x�g��}��`9��j;�΋��F;�إ���(c蛏L���T���.[0�J6�i�Xl"|Q��Oq�[�r�iG��V���N��g�lrE؄�|�Ȯy�+R��f����CU���k�����T׺4~�Y����p_���~�Bnij>��pz�Jg��n5!]�8w�{�@H�H#��[bJ�a�w��B}���������cb�!���Ƙ�o��sѨv2�v����aԂW�� �zW�)��[Y�׆h�>�o�'n[������W���<+�� ��.�թ�eNE���?���<;���^���@��S�5ݭ|-<�jZ����������dL��(��7%F�w��>��A��3}98�[�!�b�RJ8%E���C�Ɣ��XM�ه~H�Y��w��t��az��L��jc3$�l_u�����72O��g�]�P�ZU<rE����d�v�Z���[�t-����<���~JmgE"��{�yTz<��-d�ʱ��*�� ��\Ȼ��o��\#k�6H�ސ0�^�(��W�.�����!]Ymd�Y�w]�8	�B���$6�R{�L\g�fr}���$rNx�HI0�?u�m������2��zSG0�ťd'��l��&�?��|���wL*�����^���;�'}m�l��kī�h!pD����O$�L�p����Dv�<`��/�J��Q�H�5[�}�&��z�q��4]"�q�-�8B������E<W��AJ��F*����hD�h���z��,)&�2�����;����ʚ�^�"ě���r�w���/h���aR*w���x9��X�����dRr���u�Y���d�~�:�|���ϕ"�5�3�*p�Y�؃�����	{v�Q-É8��Pvwz�Z��>! 6�7 ��$QC��B �p��� ����{� �4���lY�B[�]�F��4c|c|�k�h.:��U�,�[Eç'A��M��s����Y�8/㉛Ѹ(��KW��A/�9�S(@��bG��C�ti����t�K��&������2�3����`Y������~]�;����x��mg��M^j^��`���[�S�)�Ǵǀk&�7�����Dg"eٱ�v���5*'�C�lx��q�wޥ�� �O0^H�j��u�Ҽ{^�p��8�,�g^�A=��ܬ��PW�z��3�>�p}5"�u�`/];{�]rp�S���M-���;<�0��h���a�j��n'�d2���Q�M\�H���I�r��
r�Hؑ���A�(��C7��6����<W���b�Ej��5�ZH�E<������#�3�MH��2��F"����x�qh�"7�?7��s�*9�Q� �&œSv`�s�7�쾎���/l�ϋa� ����'���~"�xL�����>
�l�=��Y�����+O�paj�Q�A������`��I�I}���P@CYn%j]r�H��(j���*X���~O!s]S8W����1z����H�Xl�HI�k�0��d4;�Ay���}�;��O�u���6Ϝ��4s�/20d_��K*�K��\rJ�������f��"�=�L�E>���Q+��ˬ�W(���+�Bdle�o"�x���>a�\�:��slb���]���Y��aY������J$�����D�5�39�bf1h Z����
6�ҳ������U�NKk�d{�&�Е��Д�L����^��(��R��&It��7�(Av��0疥i��������N�OȘ�
�g|�g����(�g^�S'�V�����<8�N�ͰZVܬ��Y�����Q��@ֶ�:��JS�:��POi¢�+ް��|�	��'KPlf���ƫ
��n��1*�h����
tӶfj1���e�S���k@���!��RV9dv�+
#����a�:��Ԕ֦��;�Fy;Y��=
�F�CKK�6��@����#��j�f,3m�S5/���P�*3��O�O��[
(��L����D��˳�仞����ǑҦF��0�6|M�� ��}�eB˄�۟�B���R;ר}��>(jV�"HƔ�\WB�
(�H����(s�i�k`���j�E�q���A_��j��uB��$���ǋ����b�5���}�!��7�£/���͞AB��>ໟ\U��	�����������v����rz��j]N�5C;�;G��Ƹ,��f�<�Zy��N~���r[K�Z�&z�+��`��m���cj�-x��oN��k}�с�%2� �CCE���zد�!����J�$�R�^
.G�Op�wQ�Vs�]8a�&���Q�.݁(F��0<p\�7�m��{�f��5�@疜r�r_A�q������T2K�H��w�����Y4|4z�t�hP��^UQ�M��waH4|A�Yha�kyL���7JFz=����`���tO�Y����\R'%��xVU��*�L^|�~���w�����Mv�]Yo�s�c�ǀ���Aj�+�W�údz�p`C������Q�G���Uf�&�c�P��Z�V��]X���������L�/�.�OUج�Y���V��)!_�4��`=�S.Oe���K��}B	�@J�<
 º`�Q�i,m�B��g5|[��ֶ�}:�y�͖J[y!w`�z6d�8Ϙ]�ܱۓ;:^��Z�C���E�A8�Y��Vݯ�UJ4�}s7�՟�w�|4�XP�������E[勰!@%��������G6xKu<Pπ�L��X.��8�q^�V�/yr�D3/^[�^J����K:/�)���J����WJ�cČj�oP�8LiSU` 49������K�NF���B���� fH�K����\��{��� yS�V���-�>讥����D#�h�=lh5N",O\t�5��t�F�j)L[s_:N�ˤ�,�_���06-�p��5#P,�O8dw��������ӣ�g��C�lU�����g�=�0�˸�Ӌ��鞅u����jr8Y�5�#�B�w�q��=�i��J�U�y�0���Ӽ-�/�S��Ŧ���HL���d�᚟Y�
�!���'	����V��6z-�q;�O��t.�ҿ���?hъ�0����f�����$��F��kL>z%_�a�n���-��s$��kR�8�F0s5�)!�u���y[���${�rv������CPy�w�}Q$�}��	���j�9�8����P�����G�|t���+StsL��L��;�<�]k�u�$�L�xt�^��~	�;2���@R���8�H�B�l�6�
��q��6�e^��ʣ�:�]!GR
n�r�������6�0��톣��|e׸���Y@���o�Ѳ�T��w3}܄OX�[��88�����p��*|��NO���$��Ro|鲺�^ـj�v��Qp� ��}�u��Z�C�.5��7y>���f铁����D@h�T����eX/��y�}:��OM� �,���Lq��ǽ�+ake�Bz[�|��wĔv�KA�н�?�~u��U�)�~������A'�f����tY�z��<O���/� 0��V/�qũ*\��O��M�S'�F��_~�A���4ܐ�\Nr��ڭRײm��P��	�f�����;�8�9�-�\�岁�ޗ��z������.9�8���$��4;��������d�6�hO�`[��̭EA�e J�y�u�Ü,O��N`��֦:*˘�	vʻT������:���{ h0p��C�<X�"l�p�rքoU��������K�)�SP�v�wV�g,Tf�JN����tj�d��m>a��PLR�^��L�ቈ#������>~�G�}�����g;wd�D����g]f蹴��Z��,u$ڮb�D�+3uu����:���q{�${��-�P{�4Q2����lݘ�|)�g�'���K��Q£�w	���|�=��" �S֢���Qb:%�5��]ܺ J��9+b��*�؝��l*��k�yZǶv���ΰ.A�*�7IEW���b�(�_�m��CK�L�q{X�(����E��v��li�'/��j��X���pC��Ρ.f�I~ׄ#�#��>��Y�����̼��Ț>��Ȍ"+q E�0T���re::�L^ԧ+Run8b��yV��h��c�Z��e��{��S��e{�=Z�?�eN���y�:qo�ҹ�(D{T��4�{�e���n�%q^Z�DW�yZ0\d���S�;���[�h�}t�o;@��5v�.u�g��9�Z�\Q�=x����,t�d���lQY�^hnIc���i�QM#lE�˴n�.��+s�/� ��J�Et��#�`�7L�X�}��T[�|�����|�G����߲���|��@'��{�Y�������R��������
�,�7"�j�
�d0�D��������G��h��Qj?�ޯ���U�[R-EH��I�aw������du-�9���z5]��yx���͜���W�}�T��Ɇ�B�/l�E$�
�	``�" O>�cc �h�kr�lT��c $D`�1�Ԃ{�^Ĉ�k����& �I��b���6��,3⫿վ��X����%���_��GFYo�[�ZeV4�q��[(�Z�L���ar3��B�+�@��*wo~����:���� Z"H��^6��$���В�x�Nƴu�� v9���;בNJ�;l@V�F�$�Se�,���ߒߎ�������겔t��/\6R~j�o���Rġ�C��=����K78>]������<��Y�Œ����0i�D��W�MAp���U�;@L�T�����T|�E0#�W�C�������cG�"�΁DM���9��B#q(Oַ�HR��.�32�ՔfO�Y�E
���΁�(>�UhU���@� � ���,a�yo�p�m[�$�X�&�
�V�b�A�`A
{Y=�jk(�5d��4,�����>S+@�7x�O�mZ�S]4�F K[�Dϩxפ��V?Ok�)v��NmE6�����@7���*�1�8@�zE�����O��
K�/��"�ȇ��_���V�
�ل���Uc��������]���o?Su���d+����(��>
�z�����L�{'i:�3?F�w>�xN�ݲ��%�0�2�� 5��<C���K�j4)�/�dݿ)���b�]�rb�Z�n܄�ڗ�v�B,�cm�<�[�}_�� �	ǏEK���X����QyfC����V���(=K8q���:V)\Wd	�*�į�|,}Y?�R���?m�{Pߢ�K8K?�)���k���ϟ��ueE��O��i�����sX�%�W�6��1/JO�dO��H�_��)�0iÂ+���~�6)ҍ��������\������mxP{%��%)��=E���".F?͒If����h��b:��S}�;�9��"���W���v����WxA�h^�˪Z���ݡv	nI>�g]D�]��;Ϛʶ,�c�#.��X�׼֗�pҊ�hr�s}�`�nJ����� ���⌝ G$5���9��2SʆC�_���J48��*�Y���~�f2���.��̰{]b!-wF��Z�hvU�K�ί�G�pS���B�Sz����	����#���æ�!R� ,w����������]�(��_{��Ɖf���w��^��T���A����rk�E�(�Vr�\���7��R�P���ԷS���;�W��O��7b���in9>���(t���9+���MI�oZ- T����g�x#OF8�WWN� �&C�k����%Ng|��0,<g�o��pfɓ������O�k��';��AT��a4y��(���/@G�{o�&m϶����?�e�BQ��H��+SD�I�n�Ŧ:,���V���Q��/�w�ݗF=�l��L�,���]�SB�S����d�����ū�r�O+Q�������^$���e8�5vX��w�|�|�V�3驭94nOm��y
`vh.*�ٖ���"[��#����'��F�DI_�n�t���m�ʜ[7�I^u��E�5,�:~B����(�������Ӧ�s��Q�%�rG7XsTh����Q���]gC�Wi�hn�6Y���~��M�����4}�l��p9��ǕW��|�[[����P����lW�S��	5F�󋶜�e\B�Y
��	�^~�bF�@^�w�d���AV`���W7�_U��_K�D���"�z���(�O�ϥ� �C��d�X��:oSeb��C�tへT�)d-g!�&���VClA����W��N��(�&�z^�<v�Mܦl�?��U�T���r�ۊ���d�Y��;,F��E�.n�eى�RJ��&<F&$ޜ�� �uˀ,O�D3��(�{��z(�F�?5��m�ɠ��>�uЫ�\��(d2x��d���W ����u�����{��/�J��9�E�;C��lV��,��{�4��g�����B*��(��Y�v�&��:?��܄�6�d�@�gXB�j=�węB8O.�:T)>��1I�|t����m~ZAt�o��@��c1Ѿ��r��(��[�'F� ʳ̐hj��8��1�D��(}ݵP!���� Jp��iv"|��"���p����q�������Tms�:���W�,I/e�¿3�۝�+���Xw�6�pP�2��7w�I�;������s�����_�G��z�_�~�c�C��,�h�۱�^����oC�@��W%��y�qf�Ztid��ک�h!<X���(%��X���\X�/׎b��D��V������.�	q�B��ݞ�u�<,H_֞�3����n�Gd�?�4VBC�B�^/�3�pW=���2��J��z�� �y7����ҝ�Ms?U�V6q����/RV�vE�s�E$���.r��<��(����&��F���a��GM�f�[z�Z<\0����Ɯna��5L�m��zs6w���S4�I��?'#(-xE�/�X
