��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s�����נp�(K�n=�̹v�:X۽�E��l��A�	;&[���f'�#�=0��C�8'if;�3!��_42:��*uP��G�zx�7pXz�>̹�eX]��9:\rp��r)����84E�)�X��"[��l��,"Y'=�
����V��X���;�z:���"m����_�Q�k�Xl��	�S�D���ː^��1X�����T�_+��#�
;�KYv�J�����qv���O�MUa``�y�:��b����qo(g�#�D|��+��o��y@��^4��6-a��e��Pe�\OiJ�;g��5!߷���zN�2�/ //��PF��hc�����v����n��G��	tQ�u��`BP����Sjcb"��.6ù�<�hD��� h,n�{��|T#�b�	��`�;�=��o��?8�W3���X�an#���ǤY�Vg�!nD�1�_�N�����-	"@	�1�Qop��I�Vw�5�{��� n��}��B�z=�F�)���<:��͉P��&�^oO�!�#)4%�2��L�)N��w����^���ta/z,��~rL^^�h���\oH/�N8o�%��cf5������LLRC�+��p|4ܚ.�It��F�{S�2�z̃���4_�-�7_��vݣ��!b�"o�5�;C�ul��SR�8� ��@-�Ԟzd�olEO:��{�-}��u���t�7���P�`�Q�$�Ś�w�X��>Y�GU���F�	;:���I[ oN���I�p�:�s�a�}�"I5 �_�{x�j���U��-�2�/��F439��H��ZZ��FDrh�eP͂��{���@�f�胚���^EZSlt9
&�/N����κ[X_���.�%Hm�,'��B�@�#��jl����Z�����(|�GM�{�?'þ�q�%��)��"�tܑ!O��0�! �5�6�����_HtgOWX�����>��m��=T�b�>\:i�y�y���Q��Mc���)>��,N6*�x��]�Z�L�)�Il�ja,�VR{4Zr���֎u%X��^�![�h?C&�z�$�y�S*����2K�-ˍh�_#��,�p:$�4^�J��<�u� 9`��ԁ&My�T���]���^��gL&(���'I���!��wE��L][�L����?����9�������M�+���TV؃�A4�F��v1����.��-�����:��v��1FeDs(R�V��
M�?|�S�7)�S�Sџ{!C�̺f6�W99��Ϸ�ȷ,&k.��M� E��I��<���,5�I�ȿ�5�������M�^��Hl�=O�^|�9�7���9�$�p�m���
˶p���ܹ)y@\>$kΒ�E����<�&e2���pEO���C�E#�;�2��|NV(ϒ�RSoC�q�	�G���x�I1n��}���/G�a��[Q6��g�9#v�����ߪ���葟VU�<>#7!����>M�bN��dāJ{���*@��� �=��Nɼ�_&��3��`E���=�����4�~����Rm��f�����`�M�K��~x �$]��H직��I���M��Ƶ�Sc�B\�S����>��M2T�x���,3Jܘ�Z~�?P���+����{.��A�_q~����r`��:��l��a�$<vP��V`���o���3 .�?��<��| �{F�p�|�y�5�7�`���>�)gKhW�:k���hg;�]	[�͎�<���+� ��n�(�Wk�q��?�����Es片���^AZ����(><� ���C}.i��6��w�m��B�LY��|&��PAdO�c_bB�J$�� <�e E9qh�	�́�yA�B�l�Bք��6#J�s-�5`��ӑ��a��Lx�Rs
:��L؉#.^�����w����8�9w�Z��QU�Y����4\�=���Y��<�⌑�$[��6b};i �?.,K+�5����<˫��eģ|R���Uΐ����7��y�֪ KDeL��[p����BL�FN�����#�� ͋GbD��m43�Q���ꂉ�(vi��Ј���Y��+t��td�����&9��o�2��<����(��4Ǽ{�Gw?�̹����,��ڃ�	9�nD:=�@]�0���=q1`��m۔���́�P�!F	QI�%��s�ߖ]��*��7�,i�_�9�l�P���|��UZ�2�#%�h������3��~�c���m�Un�/4����'�N�H�;U�q���N��cPqԚ�,�ѳ!��M�:��`*_>������
�Uj����������@�i��5ݏ޴�mF
!�����P��N�:BN����d����UC�iH��$@p�ʠ�Jl���7ɽp���:��f�(y��B�	��@m������k��՛���%��D��iX����+LO[FQ�Q}Ļ��ơ�-rc�.���2�)�ݑ�1�iKa�P��i�<�q����.�(���X�����]�"����e�~��T 1�B �@>O�i7u��4�ϴG�-C�Fu�n�:��3~ ����d�!�+���@i*�~t���m�XS!r	�	A�B�o�����_=��i�sHԌ�'�w�x��_a�����u˗`Ut�"���I����@_��&�(��R��A��H쬔Eퟟ��1X�y�Q��f6��L�Kl�6D?��Kd�ǈ���<��S���D���eQ��A=����1�ʈ�TG�%u�n���=�;/������&���4�02��X}V�s�Zڡ���)��쏇w�̭.�WAvD�m�h���i�-��q��nϥ1B�z������BR��2��B�=�M�	���?C�ȃ,�׃�R�K������	���j��N�1>���>�$͐��}8��T������WuF���蕭91��Ƽ8�Craת.�.�@<�����Ӕ���+����IRb*b�ɵ�����J�_��j�|�e,�A�:~�����<8�_$���*h�^}�v����ȅ��9�Es��s؀�Æ�g@K)<����r���ຒ�:���?�?�5��n[ī��QX��g,�}��@{֋�v%�ے>��A��R�+=�,o�5�?^R#�L�����W0�R�1����#�Vz&�%�Ʀ�c	��=�E�uw"Vs$S�-׮�ha�Z�4b�,Eg9g��,QY�v�I�sn�j��*�H����iL��&�r<t�7�y���F�,�^�l "��;��7&�G�H�BɎܜ�[�9fz��j� �b�tr�	|I@ٜ§��i�P�uMv�-��r�3"��,�)�����]��E���4��XxXv�U��L���0��CjT�jV#�o4���5���3$ �X�����i�@m�?���:����)=�h0A։��9PJ&�tXq��Z�2'«��<�!/���@]��V= x$�U��pӑ����k��tM,f���]*SeɃb�n�J5�����@�S�=�D�Q�Sᰡ�#X7F�a�y|�����=�O!��г��m�_cM񭧮H$�I9���+?0ŚJ�;�����N� T�<����c`���Fa�z���dJ9�$���1��o%1��Y"���9��1��R��$�3��\��� **`�B�Nn��&��4 �^���\�g>�K����Ɵhg��Y��sr#�g�r�@zl<���^�_X W��5TݤET��uG�^
����ٜ�1ڞe��4�'���R�T�{2��L�e��u��$�zNbmA�R%��;OSٝD��cSM�t�.V��Z� ��'��i�d��al�'S]��h�t��\,����i@�V�Qc߂$�O�nE�m����Zf�K#&�{��s� w��J�v�7�ӣŘ�$�Ꮥ�[�_�#8R�5�k�C��Q��H�Q��g���B��	[ ᠈ӅB�p�x�V�_W=T�x�:�7��9�b�K��� �:�-O�N <�j�q&�Zf|k�a��m�	�[������;5>b�:��S�����P6�f����f��?0qo=�L�_�6D/��󊰀���*�|7ùfi4w{����w�L����eTw��"~��]����"�+�θ��ӄn���H6}6�R�D1bC��SQr����]�����킧�(�/R�������\-Ӹ1�Q�1us�������O�bx����I��9�,���Y��b���=��RA��ɣ�vT�R�vu��L�]e��Q�Qu�xY�AL��oz�B9*<�Ȑ=�72K�� �	ś���%�CYu��@"�,�
qp��hTQH��^���&��'	/��tL�l6�:�)-�T�嚄��K׸�n�2~O�'� Z�3Ba	�P)(���T��e����|3��qX�T�)�ҟ����-�ES���'��j�1��`������d"��	X�g�b΀΅�k���yGh�[G���G��AW���,ꑱex��Q}vu�9��ɱ�h2�yF�U����Tf<��ɧWo$�W�� �t���aA���ڎ��Q�H\0��ܹ�˸V���]Y_.@Y@مZj�$#5���'�~
�>����x?#�K����P�d1�ʪ�iy�mCK� ��ۄSom����;-��:'�س�d��n�A�i�.�B>��@J�QT�j��D��*ȕӚ��|){%�/I��s�F��['6�M�'����O��|K䰷F�D"��Y�=H����5�I������@�^�3��:�`��JT��!��j6���k���V�gq�WiO���<�kɦ&�x�<�v��P����?��9O�'� �����e�4?�uy?�PW��Mт�S��T��\�����=!�g��q��M;<I����){�`�Y%R�l�X��:^)N!J�{_2���җ��'
j���M�1%Cq��4��Jԛ��6��y:v�s�v{��t@��!�Y�	�î�Gq�j�m���C;z>�U;VthKd ���'If-q$"��5`�?�7�0���F���D~������LQ� wE�-lc'��>�<!���Ŗ����1J�Y%u���UF��<�j8Il�]Xq���u��2���Z�!��-��:VJj��XZ�c� ��za��	XY�#AVq>|�Kr�����?��i%�ה��h��7k�G�c�5��֡jyK;U
�Ϳ���o)��Y��;�ѣx��{�~��XR/[�B@{��_2�hdd���i,w(Z�'c^ز�Jg��1��ǚ�=�u�������Y�sc8S���P�0��p!����,�y�(������}�*uX��Z�[�����`+�tE�|Pwt4n�Je5Le�L�L�dB��Vt�E!s`~��E�e�����Z,�W��!�	�bԮꜧB���E�Ut$X$\�X#
