��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU����ax���Q����.�Ā��{�&Z+�+DZsl���Eg�}��e�č�%.��R�3���x���S[|fVs��y���'�>',�}��nXcx��Z(��8nmX(�����!%ˇ�T9�lF�	��j^lU\��H�չ���6�p=īx�H����;2�����tN����Īr�v�>�_�dC�coG�zp��q4��*��Kh���xR�Z�vI�G����K(֑g8=��#�(�5XXU7iyΜ	����$O���0�j����6��9�J���7|�64]1LC"����P��\������~'톓���L�ѢW6� }���ˬjO�Bbp��VY���D�����&=�{�>���U�n`L8ah�0�MН�N9FdF�������g(ӌ
xy��	����sW�d���a��3+�K2��F�V���?�_7�4U	�~J��7���YV�U�@����o��Hص�FĘ�a�ΆE��]w�=��Jl�~�T�x���M����,�����V�>�X'��Y��8U��x���|��%��
6&}0ʖ�"���D����7�D�u@�����a�0�M��T�z6�_���N`#�i�z"^���cޙ�7(�f���x9��m	��&E �V?4<�X ���ՆZ�j�S.�y"����~�"��cG;w��q��i���J8JǗ:�2ȏ�&D��p�F��O�w!:\Pu����nX��`�9�#@�j���'礬r���QJ^��yE������l�V:�~ �ٚ����.�[l�F��誙OO�W�~����B4ӻq��<���{�u/��!W���l��4���8!�`��ܲ{�5��v2'�ٖS3��-C��!�j�0QX����Mv\~�
��1ی���
����Tm\��	`@�Gk�u|P�����^�)�):G��. ���94��J��
F�-M��H Y%��ߔ\��>�V�-㏳I���{~8A���߇�.ƭ>�?*]���-N���;<P_�XQa�%�_��9>���#i���H�6Q���2�{��	8�ø��pZ!&���r����Z�������[�M6��J� .Z��L4;�h��_7�6Hl��&�״@ɘe�i>��OwW�m�3ǆ2�Bl���8�Ҩ�i0�OGTX[��y� ��}%�2�~���ʦ�?��V�J�쎛�@�X[x�E��W�	�FdsP2@��w�cX�$ڒ�X�"NV�xJ�(+��P] � K��]'�ﶍtO }���Y���hN��ˌ���Q3�s6�@�z���9W�B���Bq�)K�i���3��I��_m�6xXe��Ϋ \�Nںm��T�!S��\����{��7�*,�)KOi���]/��rw�\��2mî0��w�TݔD���v�2��l�Ж]#�O2�Z���E�գ>�����fg��5�G�����_.�7�w�F�a�9���n/��C2�cǩ�����#���5��툫����O���O#�����G�wEԂ�%	<U+�(	}J�H4��}�z�T٬�����,*>��[�e��][��\3'ת22���q��
���I"�B�M��r�V~7i8�sb�j_��J����A�҉W���(���X�2�
��5�1��S�<����^V���*�z�ea:�
�[WΘ�T���R���)gj"	�o��>{��g���@�87�� �.��N��JV����c��S.�<���3d�������TIg/��g��ۈ���}\<"���¨��V�����p Qa���S4����SFl�O�8$�O�se��f��]��w�Ek�Ƿ�����4V�.��Ħ��x���S��:c��I�0Βd�~������D��z,��{UI)�Y�90��W=L<
�L�)$�lrL����i\xт�u��ʅ�>�v�mm|ĳܡ^tY�Nl�y,�I?-PD��|.Bg��r�v\���2@���ÍA��8��h�I/h�7��:'d�>�*m,�ێqw��r�k~��O<����M��J@ͬT�-l�a��f|2ƍ+���m�T7��?�3gi��F��d��Ho�k"։dETe� ����_�"/���LKEPK$� _cN�r���O�	���E��S$�c.d�h���u��mK���Tm����T�Q\�w@e�Y��~/�2Q�ZpT�ѹ�d� C{��XB����s!v�W�!�9���:C���`��=���-.n��Z)�v}��Ɲ<Է�j�q�C4�|&Oဩ;)���˚��$�-�CݧI�
G���+@@}����d8��]�T�ku��2M���b^���'�x3G�?��tO�;���B��b�ǐ?U�&��E8���V�@-�SJR�։����]��G,Y=i�ݎ�IfL
�A,���=��<�eY�Hn�N)վ9���h���v1��)�'��J'9�h��k]Kf���zF�
{_��@.}������g7ۊ�
6M\ن G�*�U��6l�bf_8�B\~��j$=��Xs��G�M��v6h��C�}f�{�h=n0�	���YP�ퟓGFَ)vO��U�)�=�Jzk�R����L� ����	k,(J��W?� �Hw^����eFu��[�Ō��sb��(��zl%����f��S����o=ӭ\�>%΃%�����fnIF�b͈26ᔆQ��9aW&���Њ��<�z�堿��j�خ��_�B:�t��첃W�&/!g	����2�2���I�_�2������*l���kJT?@��L�,E}�!{F4��d��Ra�Ԣ�z&������g�mZ�
<c�%�f��9)���96�O \t��w��@D���|�E�{8>��x33�R��h��l��.2�����0�>�q�a&�K��Xr:^2Usn���k��~�BL%�s]۪�wۖ���O���G<�$aWװǍH�:��U۟�e����?2�4w! �%�Hv\9����_2_j���#�c�1j"|�e�'�#�Pd�E����:e�����s3����t���7�voR�$O)Qr�y�oY�`B���">H̠��f(��l�Y�d�#p��G(dm�!�zg��z�"���O�����C0�v8����tⓊ�a�D�_����::��-�J1���(�����e�pP�d)u��-�� ���E�*[P�j�o��)v��OYk6����ğ�	m��V 7�Ml�󔄇Ƥ\�vR��ü�l�^�`F�F�feS)#G<�6Q+�X�?��f��L� ��L;Gm/0tf�E��9U����U�u�������,���j�G�44���(m�ߎs ��;F�@��>gXn�ֻR,Dv?ڝԺm�K�?޴z�P�,��Q�H�$�5P`�S1�H�M�h�P^F�Hg�O�k^A��OX���2e%aV�щ�g���0W��#���{K� #0���3?	d�S�ð(!�Q��T"9W:��3V�_�PY�'�Z�KXb�1���XA�}��V�t�`7ʿF�E����dOU2P��b���q��;�X�V�p�m��Q��;Y�B�o�M<��p��n�n_�~v�۶���b������h1��ÿ5��#�Hb$ןާ�,*e�, �&;t��$�m��U
��9&?<z|� �A��c�f��dZ��� e��Ĩ���3ftX\�$Z��!FmP��9 NclsRQq~�!�n�f-�a����hv`��+C"Ӱv	aͼD�)ѝG!���>ċ������<2��h�c��,�t9)�aM/0&�:y<�������(?%m���CU�}��Mb;��O���^�G�a�IŦb�%D�Ya��!��6=�MR�,�o�g����f w:A6Hy�*�4Q�����Y�~4�mI�$����@)�A��&�`��u��f�����W��C�+V�>�li������B�!a(����5���D��I�J�!`�����
OZ��}�uw
�Z)Wf���:,T����1-a�0��P)d<���-��ԀC���ם/�j���Z���L��9�W�V=���'�-4�ԭxE6!%���^齱k��|xor�.+K8q�����||�#�E��̉��b�n#���l ���҆��-Ԯ��:Ӽ���|��8��-Wof��a8B��wI<���-�x��$��`���T�~�'�d�
p�> �1�8v���j��tz�i��
~8-�0m���H�3�#ܶ��T�q/���^[At�U&�2�9p6��J)��:��_��3����]�5�Վaqg�ы�ZQt�UZ��3]9���q�i�����^o����u���Ͽ-�ez�#�4'�	�,+���8�|�v>O^eY.��YF�o��%��1�Ǖ�{�嶄�okx��M:���ʸ�;F �8��R���{�6%-�q�Qj�K��+xd�;��~�ob4��x���ɿ(,�b}2�7����~Ӊ��������-�<�(eM�K��������:��>�l�*��TṳM�a%�\zh~��(ȳ�L���iD�h����V��gX���	�N�ϲ��.���5��K�pBi��(Pi%����`���:j_�ڱ�@۱�j�6��ջDD �i#�X�S�>�>�@�:9ڧ7#B�Z����DB�r���>a������1�a���y�	�uʏB��(����.�F6p���s(��I�}	�J�{O�����`%�g��B�$��K�����������fA|�3��o;�9����+�t��]//0��<4�E�]k�����v�QV3d�\�Z��(�gJ�yp�xWq�o�Í䁏�I���LP�)�n��7XZ%cy�i�I�r��.6'7%;��H�:|:xU�;ʂ���y���c8^F)�*�N&�b��e����4�r� �*n�
`+�w1ј�sODh���bG��ݢ<�,(q=�^/-��NLP�5���>0>�X�Q�.��Ó92-�I�m���\V+TU�|��a.��'��
&[c�ma2�*>Z�vןO\=�U�t��E���=j*Pq�l#���}ozԹ��a��@h�����A��+�O����~Q+O\�<�U����V�B����>�:��Ӭ�Y���5wP�L��P�u\�
���������2�x��mo�a�l>��w���r\y���R
܈@]�#?����=��7����Rf��#q�>%�i}�s��2�`�M���u�v����Jl<��c+��.��|"#�z��A�(�0?����"e�2i�$����t*�f�nh����PlhA`�`L��ە�#p�Y�:�K׼!/f�0%*]	{���V;����(�':z{s�a&���/��;ֱ̻IC*��G=Ҡ�2i��U������8}��1������~�p�0Y��њ�m�dW��$��i��{����
�Vt���U��3ӯf��nr��D\�mD#B�/��XKR`O�_�G�Lr�����Y'X�Htz�E&�s3/ot�����5~�Klҍ���.f4 ��u<E�u��*�O���q��s����/X|��ʳ!�~�Iw�&
!��Y~��ګX<m+|���b&#����C�k�)>�D[犓C�VQAOg��EA$ʚ�t�Ve"l���=K����s/ @��]�C��[Ƴ�-"���	F�$��թ�hk�h؟>���5j�ݪ+g9<J�aQόd���A\�I�{"��Y�4�z���d#�\�^Nhr<��{N!�z���W]��xc�L�7�ɧ��� T�Q����^��f��vDos�ﭙ�����DȖO��ۛgB�s����Pf�ᔯfi �~X�)��@�VU���04�x8>�	�\!��A��&�iyg�&A��O��b��>�7�E.\�=RP4D����F��E�,;�"1vÝڝL������"�d�C{ss
1h;S�QK��m/��2�r�(My^	hp0�|U'k��,!�s���C��Rk���\�ZF$qL�6M�!	:���˧@����L��Zp��"���z<�2ϻP�����w��ͪ�%)|����sP!_��7�K�*N��rk�j=�G^�D�6���������@w�-yZ���{{�(�	��N5�<V�m��6��d6{|����v�9V��"Ge��A�i4Yt���E*Ꞹ����G{ZN��1�#݁ߣ�7�YF	�B��MD���0"��X�����{<��'��2YXu��&�.8�RƸ#P�R`�l6B���U`����k�0I7�Ykti��!EY���K�z��3��o�w���w)�'V�ɀ���x����M	~�SM�ig�	���9�cɧ�6Nd�'�T�(}�\Md������t��(����>���	��J�n��W.��Ű�dR�<a���Cggg-�R�8!����{� n�c��o�^@�*��;/m
ůNV�����yΆ
܄Fm|I�#xQI�W�R�y��I�>x��-g�+,��'��C{BŮ)�>�c"Bl:�E?������a�;\�N�����I.��g:��"R4{��#�\
a�]�J	T�+��y�#�Ǫ���	I�7�.���t��
�lo���7C1pH�%L���B8-`�v&�5�2�I{�3R��*v���$#� ��2��pP�SH�p�`~�m����a�����tXZ��,��i�lN2j���΢�w+�Nz���-ɑ���6��6�:U����Z�x^�Yt�R^J������z��$Cb���z�f���$�H����5�v#V��������&�*��.�r��s_��] �&k{�9t�����vu6TgIO�����CYcC��4��y��	ˀx���P0�,8�]f^��z�Ӥ��]�ܸ�py$J���jb8/U	nqJ'1�(�yB����c��It��s{�^����:��t�9��]$����YW�[�6!f*��;ơ�Inp�q����T��d�6��&�*z�:���oL�C��1��|�J$a��(؈Յ���Wu5�����wn]%l�	�>*��80>?nb�-���bNe��.��ɥ�b-��c�������]Ĳ���x�W&uԀ�t)�C��V�}�����n�n(��_L�9�v�9!��n2V����@I��v��g{�o�L�_���LD�-�z1NӢl0i�<ZI��l�͏�ZdYj�/��P�$����>]	亥�{�3�!U�\�˨L'�<֚�i��8/�rH�0�O���ܡ���(�5{�b�1�~nC�_T��q�=�jaEȾ�]��\+;೵F%�F2u}Ԍ"��ןh�h�/�4�`�\u��(q3hK'{̐7YM��&���ѝz��,(�̯� 2�N�{͖o�x��g����Ю��^�r���k��> 2Q������a�D�;V���]E=1�Nb$3�r�k�u�����C�7��o����g�K*3�,ۆ��,��>0��)��薲v�MX�A�c�Zty�.휲ZWoH�Y��(QgP]��^�#<�M�)���h�}x?��q	�T7���ʫ3FΡ�j��N���9/�ϗ���GI�8R cjH{i����{P��w�D�m��n��?�~���Ao�N���CKe��?|e	�h�M��췭fM�CkhߥX�8Ï;�K��⢪;^��ߛq�q3��R��S�tt��F�n� "��;}� ԝtk3�ɠ�GaEP�S��͞Ya$�h��G��`C;ᓇ�kL�v<GՍe�N��q��fa:���,�u��Sj�_~ꘂMlu�3	�S`�
ﻷ�"vۋ��S&n������J�(���m�c��Ź-Y�G{�U��цGy�?8q"�6�E�,��{����	������!�Be�(̑t�P��� ^(�
ը�fxu�a_8�!Z�>�����:(�6�b��m<�N}l����cCJd?h-y��Y53笼&�6$>����V���/&	��e'>1��CX��/�5s�����T64�uȑySb��Al�>����[�F�!+��q$��]�vW p:�Æ�(C��3	�%΁R!N��)X�L���b�G_�o��X��ݔ����pU�S�D��Xs�6���`��Հ��'q~�h�P�&~�)��9��%U�q��IW2�˨S�!�o%��iX�(Q{�¶B�������$�<a��aO)+0��qB�6l:�<B�����)��,�J4���Y�Q�/����p���ON&$g��nJ,�3~y7��W��W��|�ˏҽɋJ�)��͊�q�G��!цς|���S{| o|R���홶�]���FC����\�a�c/�燚p	n�H�:q��qP��}�<�R�8��i��KCs������-���-XC�k"h�q��@�G���U��ڃ�������0x{����J��SLhs�"@���;�~
��q�>^*���c�gq����(�l7qLeɒ�;��������jHN�J2����U�e{S�4;O�ňs�<P�k������=����'MC����E�2+�7g�l��t]��dfd�Z��+��z������.��a4��/S��CQ���6FnsЏ��4����Q�h�pq�민�]��C"Եcx|PK���*�E���4�����hd؆�ᾛz� ��~���~}��k>9Q������*ppH��a��s�t$�ro ���,�4{�ߟ�jX�p���kƯ��Q��������+�c|�"����|�{ q�`:����z���)&v��7X��|����r8�.������ΐڲlq]��R����k��̑�K�M 'N�Oh��.���E�vZ�d�CMId7�΁�E�dD�6�\��x��8���	�&h�U62+A��|�x���AR��,ϣ�-|`�_q(b��!��������<o�bf�zn0��{�3�ؗ��oO�:�`%�y̑?���K`�Ï���ۧ���"���K9gd���V�1HZ~c�#�%W���>JX.V����<���4THN��EҘ����v�Rv�Ķ�6��>�x��/������V}��y���J�yCH��R�<�O�sO��/�K�8�/����4��ޓ���W�m"$��_��y���x�$�aѻ�{���[Yg&��_*dO�7��/Hylh���5��ň�l#�F�%S`�@���cu~~L�2�y0%���rg��.��gS���%��?EKWҶ��#dIE��?� ��*�#We�O��@_���)���!F�����P�3��m<I�U��kR�>��N�fC�����������֘j��B�(d�>2͡���v?֞A6�̌}�����o��f��_**��d��$5|s���6!L~����n�>�ʻǦ��S�D��D|��G�bg0_/Y��"{���@�T���w*��X��{�gkT\��c�-l4� w�$� }��Y;ȫ�"8gnW�俺[<!x��O����T`�������	IG���X+�:������z���
	<��-錅\�ϒv|�cL��+Os�䞌�>Tӣ��K�ӝ��K�23�斐�y�^4�V�q+�t,U��חM��qHt�������ؔ]�98�����]	.���}LR!F�6�Ln���R����v�_;�F�>�����N��Q������g�X�Ș�Қ��}��ƔPP,S~��y��IBIN?������@�yָA��۔��)�м�q.�Z��)��"�oB F^��u,�G���>Vޔ"]��, 2HMu���]����CS�fۤ�vJ�>��{V"5#�Gs�P���=B���u�A��>xӹQ37�g��W��#�D�q$9�GB�5e¡tJ"=�^��k�����V\\�����Y81��Ǣ?,E�o���wz�*b�8�A��5�\f#���5� v7GT�F���~�"���m��?�2L���[�:B]�z{%+��7���Y�=�D�#EQ����cb��b^;�e8�5v������|��=T
��N#�Q4��	�O�ꨓ��bo���4b[N<���Ș�Z��ܑF\Q���!�
���k��[���ڂfm �¤a���W�\k�Z߸ey�kǶ	�wUQ��:,��-g ݼl�ȍ#2�	�t� ����H���g=��`�v���7�Ш܁�ʎ6a���-��ά?�'&L>����i���/:��Z{��~U��:�������-�|3T�~2�o�O�F�c��8l*�i1zk�2TR�%	��"!����dc�q�D�\�>�`�OӇ��HR.i�>�:���3Gy<<���>�z�}����`�����B<����Zt�	��TIx�}��oGi���v>�d`+?��d�ĩ(͠7\VW�G>2?�o�C���i@ӡ��'�/i�������������*=a�r����������V���=;�T�f��g��,��볯B��CoB��
��ܯ�7��r[�����JJ����oS�sz�:�2q� ���J��2�� �q��v�ʰ��^��3*Q�G?0��z��o���%f��mx)��Gä�����Q4�`JL"wl5�)ZW����#+�\�.Yi�*��2k���~.����+=�C-���V�����L���o�E�	F4ھ�f�1�d4����[�o�?��Z�[�G�/(���F#Ewf��aǦ���B�܀�w�5i[:X�M�VB��*���9��"S���z�kE8eBE�up����e'����ط͸���TkK;V��X�[b�㬥��ϭ
1�y������'�����'�M�άH����(�	�]J�ɴ̹K�N=�������U�<D�!�.吟P��f�aK�G�i�
)�QOR�x���;�E������|~�����d��]iqcn�9
�?1j�P����M�	������U[Xʀi�2�kU$��r�{�$(}\ tM��ԍ�N���� �����JλS��#�w�V��ze$si\���/.i�J�OD*e(���c���|ދ�GOSٍ��J��4�ظZ�� ?y��I_tP���X8v�J��i!�xe39vR�1#T5�9v�H.����j-�.���9�V�7�V0��uu6�4D	���A��VI4FYRO3��1��q �Y%���ry-����T���ޘ%�Ïu��X�nq'ɺ��pѩP�(a�������S��>��M�e��]�4��:����(�ą]�i�ܡ�OϺ2��u����VA5L�5��R�T�8�˲�#Z�����p>Y���[�M�O�MMj�q�ښGG�vPS�=(�{�q�ͪm�5��d#�"Z
�����2���|�A��CiIV3�����f�05��x��jI���A���w�ԛTd<�A����DI�'�9�!vM��9 �5ÓAơ�X_��M����c�O,���7�^�#��,��,����~o}�8O��6�!C�@nnI�՞�b4Xg�U���)@q��arΞ3UBm2�_ف��~c�v2چ�}����85$��R����{e��W�x":�z���Xp?��vjX؁��^��Њ{W6dWŘ���� �����<�^vlj�8ɿsB��>X�����W\ ��e�qa��l�d��Ɣ���^��>��P\\<IT�^�R��YS��ϙ+ڃ�y#�����,��M��Z�9�.�����}���V��r��<+Ω)����	���~,BWrlpXh�����}�w��Y
�O�T�	S����������k~�=
��N��q��$��>��l��ߑN6��1�Lh�يw�1��1E��A宕�$�w����@X�\�3���Rl��P�?��}�p�E��SL`Qe��q?��pc�
�vy��!���ӣ	[���ts��~[Y�3�'�(��P�Y8�j����:�x�c$��+6�w��M{Y���/9�{�(�Aɶ���;"�щ3���(���;L�a�������Q� ����{�:f	�+v�����u;D>ݺ�6sXӵ�Z��cB|�~Q�������I���$T�.Nq�m9E;���v2�|����%|�F�}x~�^t=����Y������f��x�)䮆
M�:>�e�3tƥ6�cm�c5!�f�g㭼�T^=�ش�d��w�=>�����>:O��P[O�K�g
�pS�Qʯ�Z �;si|/���qO��O+����Ah�D�`O,�7t���C�V�a�p�d��^��.K��8QY"[ӛ��U7ӽ��[�J�j�Э�Z�#W���Ɋ�h��L:mܐ�k��	����zhS��'�i�6Egu2*��WyAN�~<W�c����}�.��<�W�F� 
�;�伖���%SG� �L��b/=�{��?J���$Ŷ����s�p!����a�H�װ|x��6rĨ�����-	�]�=�M�!G;�kB�lq�$�:$,�I���(�rF��zY��S5�J�v	{�t�/�&p1S$���&A9+?I��0�b��tŎ�:F'Va>���.-7v���:��QO�z��O���+Y׸Nr"E�^ˍh1%ku��0��(���w"���l0��O�f�[u,��\۰}�8�]�i?}�����|��!��o ��6#{���{S����n��T�JRm G��_佲+��J0)����&��{�5#�QG��D�]V��s]d�.b��3��!OGu˦���^?<$�窧���n	h��8��r�L�ڇrҭ%���ל[Y�V��j��������T��*�R�[?5_��&��M���	V��nI�Q��g���b2���!�ӋH��1 B�ԭn���y�u:�B��x
"T�����l��$�L��z�r^'"���Czw&�\�
���\�/�D-�u��#�o�%9l�?�o��j�6�"U"���%G� ,�-�{J�ƔN��8�ʘ���9.ib:�$x��<�=ss>��y�D�8r*q-
�f'����wS$���SDS�C���yO��]��`��;YS�f=�.�M��u��P���J�iU!��ƴPD^����#B�_�(¶튁e ��L����`�]�F��yHH~ ~�
e3��H����nS�'�;��3}2����Y�4|>0m�i���7<��1,%%"�{k�j^�G{�b6 ��o�>U�R3�o���,���AR��f��ߏ�x[��̆�9=!�@���g�/B�0c�|�	S�>l�	�����>�x������N�����UT���c��/�G�}6�S=$���*�奣�/�Dy�v�<��r_�ҢV}1�qb�S��*EӺ5��� ���)����,�k��5���b��#W'�3뤱�p�>�������v�ʷ����q|J�l'��K����Wo�ʁ���!E�^�%��iodlb�pwZ/�����p	��qEp\�XMy�V�M)u�Mi�,'U��a�6Ӻ�u�rt��}>K�,�S�ke����f���K'u��=����qW��Y�O.>Ā1��=�4)j�^?���R��8ar��tK[�l���ۏ�s��(A�Q�C��N4��"����ݲ��\7k։*vx�u�D��4��8���\#U�F���NQJ��!v���I�.T�����[HU�y<�.Z�����G���ZI��`� ���H�q��d��X	f* i#���AE]-Z�b_S�lH �;(��Ҙ|��陾P=��^��,[�_�s2F�+��F	�n�~#4��F*N�ȵ6%�A`�����Wly���K�I2K:��9�Oc�R�^��@Uޖ�DK��r���[^h��,���ذ��lJ�<)�"�p%F�fz�8�[ʋUʁG�=6T/<FEf��D���߀X�G0m�r�u�!��0X��h����?#���Qv�/�j�p?�5���4�(E�d�ȺBw�2�)�,�l�,��FcZ��@u�����|T2p`��U\2)��C�KI��B{,p�c5X��A�T.-���Zކ�&wɒr��E�jfQi��'DF�P�����IB\��%��0��q&h��W��� ���k���O��FX���#�u��L�S7�ei+r~J'�zᚕ�gq��N LP /;Va'�=]Y��a~�-�۾Cå����u��@L�{� M�����c?VlH���Mg�b���S]�^���1e�叅�B���gY�+Q��M�M}�%'L�&&���x����av���&�oC�d�
���-۳�k�z��d�:=�x��4�Y�"��ͼ����4}� ZͲŪ|����kZwƹ�:�z	�B��j#��E�ܦ^���0�]���*�v>Ҝ_���?����Q>y��:�D��x�9T^؈5̷�h1��%��I�"��Nsb�',�?�9՛Ȣ���`�q��]�wg[L���:P�P�$!}t�l�^��藍ۻ2h�xQ��	H���
L�dI!f��ƵR����ff|
�I�@�os����5R����&.yAx�Z�p��g�����Owk�v
��6�ԙ�U����`A�_K/kf�V甡�,��ϟ|
.��{@mi������9���?NO���3�8���z�?�"�� �\�C���"	���i˻f�1?���l	�g�ŵ�'bT>�ﷴ�_��h��.�I �����6���y�q��X��\�{F����_J�4�^�|�{��h�v����/��^XSX��PºM�߸q"Oe��h<(�=Dy��LC�֬�0������� �d�w��\�*�4@��A�?35�X�v�&�^,s$��p�d�R%>���%d��Y��p�1��f�������n0���=7�ɪ:l�tʾ������t�7�k� �YS�=Ų�밭��l���sA[$�2�Ô�F4^��`4Rפ=�GK_D��0���E��{1dc����!���@f�K]�F8<fF�>oxٌapwfԪuW��_Z@�q���DN��UhuP��=�ފd��GF+U�4*'�����l[s��a_-g�t��p%��ǅ�JǑ������#j���rͰ&�EDw��}�N3�l�?�3�j["|WT�w>}Қ�?�Ūg�#��d�d��;���$H�4��>�i��S�!?oR9�R"2��3x���������v�~�+l
�x���H�d��r\���1I|xԧ������:�i��Z�t:u�=q��^"6���A�=��U^�WІ[т�?^*gh���z����Q�P����,����(:��FV���AO[܋X)7��G�gLX�f� �q��w���Ki�q�w��$�bZ�s��mGJ��(}�gn�(�}�6DO��;�WH��6��2�G��CW�ߪN0˱��YEג/?�F�4�Y�ݍ����~���)��M]p��4���š��\��uϗ � E@*���G-o�i������N�JSw>ky;��KV�V~N[T�O��wA�,�� ���Hf^�tGFa0�&�hG��G�u�FlM�A�8�f6hR4/�#�!�D��#�b~bF�{ut���Y��p��x��������k$I�PD�I����*AT���gS|��H,��J0麆�rhF�S�E�t�q���U�.�RU��Tn[y��ݢ���X"a�~�$d���6���N��X[���3c����>�GL�g*cb��X��z��1?#��{�=Jײ�w	�˄iU���0/�D�h�I_������#�����B����0�g1fP4����KCJؑz^m��p�t	t��C�-�	��$L-��g�N�-=���Q��`��T��G='����@c�Rx����� ����t�#���M�,���`�ȏ�l�1f�~�I�*ztD,�˔5� Ie���A��a�VV����;������H}/c�8���B[�o���e�f�5�fu�|��Y�;��$�������j�ˢ���Ř�GG�ڲ�A^-0�nZ���.�ž�I���&\h��Ř$�O�$�{v�TeY��j0��% ���}4~��KfP�Ł���(����ϰ]%�B��{��&�i܎F�e����a�) �W�-�z���
�tJ�x[}�X�g�lT���բ$	��T�#Mw�q]��Jj!�ԯ��Q>{Sq`��4���\�2-�Gxu7|U��,�F��c�y���y�D�}�&���Wj�;2I��~+� �2��@�!���:Y�;`�:L=2�D�F@S/4��T9m�ϸr��l����$-(�����3��_ʵ�.A'f`W캖�f��u����d&��.�c����c�����2���Ⱥ|66=|7BN���q{�D����#�@lI�>�g]/�r����*o�t��E�y$0�0�vC�N��5�B���3t+T�<��/���\~48;��S_��w�b��TWP��߮�Y��c�Fθ�י�������[G{�!U�ILkd��#�d����es�<*g�[�:�V��zG�f�U���)�i`�� �΁_g�F��Ta�z�������u�yL`�IdA[�L�ԓRE�������}���P��2ɈQ�s�y?51���bFwv��RP�fi��P����}@���;� b��&M�ި�<j�k���<�����~��t֧!�`����_�4L��(�EF�.ދ'�o�d��T�\�l~Q]��W�����L�Ѷ����d;��ெE�����&r�?Ӯ���r%����U1��jS��3���*�۱��<�o͹��@��P�y1O�ye�"���ۙ��T��!�W���b��q�WQk�]/6���7��f�JLn���0�-��^�3s0���JuJ��q�,Gk��l5f�iI2��9n��k�����:���3'��������ʒ�o>e�Ӧ�9�;x��6�Nk5����]N��{DK��s�� �����B
u�A�� �� ��@ߡ�ѭ� ����@�P�y7%�X-pn��q�B�(b^��Z�(�������`r��獹�4��jGt���m	ȶ��1����+�9�N܃`e�/S_�-Ua��s�}o�.�ifz�/���h�Ể;<U3���,'�����(�ή��d�Rٻ��N����\Í�"J}js��쁡0�Y��0�f۩�?0���4m9��,��4r���+R��/U�����o�Ae�%������q(��LG�g��gl=��*&���٢�SA���U7"{k�$a�w���,[�K[�B�%���J����Ks�	x'�,�<�1��@��%��L�R���Q�y�"��T\/R_��^h���#�������!�RE�L����c[�\�KĘ��$d9P������yz/�:��c�������M�85d���o�\���>%��+���C�T5=��Un&��9Kd��} D�\ ����):�s����f���wѶ!ż�Rekކ7�us��?��yv3��cj�Pv�I�f�II�2 U!�C|�v���..������+�E=�X�e��RY�OM�l,��I�2b�%`m����]D���@�+����Z�9�Z��Z��E{mF&~���ޅ�<��j;�`�l�TX-�rVe:W���*�\JO4+r�BAG��g�TG�p�C[�ץ���<��E�4�xN�y��&�U�r]��;@T@����t�;zػGR蹻���0b�%__�.O3]����2K�jR �?t�֔�_�����kf6F��Y�.��ծh<����f-I��<ɍ����;G$R.-ऋj�T��v�1�FBI��F��̚�<c���S�U�]x*ֻ����1MB�H�6J�=�Qj9P��RO�!�"�%�@������~��X�p���wn�8pa�d[yF�7���-�fo?zmz���g�D�|���#��L��$�4YaC�)�4ς�k4�]�S�%>N��`�����y,۲�6%�<�>��T  ����=���3��7�G�ꭊQ��Vu>�E;qB�qO!�!SN�����cv��a�F�X�'P^Z��Iz]@�z7 =��5�𣋍V�����I�����Vqxwx;rV�����o}�K�#�'���nU���X"�K�A�RI���\�T����8�It�������G<i�J�&_.��\��oK\�efнH�-߼�iH����Z�{��+�����k���A���8���w<
�?|�~
-��n���ґ��*������Q�'���C6;�G��/�=����ĂZ<҉Q%�M��#��������1�Yn½��C/)���Y���Ug����O-,�Ȩ��R��Ҷ�j[Y�{�j<�u�n�gիw���&��z�ϳ��/V�ApB$��t↥��n�@4��`�Kz�@�2�X��)~����i�
��z����{����i0�L#�r
�������O"�7�֒Dq�?�78v[��$���cR��ҥ���!_�k������7�]�&�����}p�1����Y�,	DC���[*����c�÷�g�hs������M+*��^�Oc>6�f'��	ױ�[r��.3�e�q�W ���1�����g���3�®4���5�YC �������q�	����+ ���R��F�Z5����dĤ
�\-���gI���<�k�iJ�\e�H�	|^�"�>���/u8Xβ�Vv�g�O\>s���6�e��6�tNF��O�O%��\l��o�[w�V��~�i-P;��GA�,��1͡}�	5z��MG��i+\y���z]�P��1wAlA�9���j�����I����qHÀ��Y�fn���@��%��� F'�j�ol�V"E��X�1􇯖n�-2��N0�TU<�1h*6�l�(G��nއ֛i�p���*��A������7�����e�X"䠸��A����.��37��op �[W��(�Ǧ|�R�G�{+�v0#��TS�Y�M}<I<Ȁ��nu1'�N�ȯ�����(�L�|�ѣٷ���)@��%=r�:�/�G7�~�]��,bb��S�Jp~*"z�/fj|�Kq@~J�w[��*�N���W�Yw���x��ƌ8���u��7�s�A�����^��b��"�J+���w5����w�$�s:�Ž�rZ0ׅ��1^�Ȍ�~p)`A���l�GB
���hҥ�G�	�g�qy	����d.Ҽkl ��1�#]:<����E8Z��IN/�D�i:�65N^�@�)�U�������E������Ǐ���/�����{�+���ζI�q�s76Y�����a�Ж�2"�qǡ0�LwѪX�C�jV̎�m�y��gf�疄�h��FVW�4��7E�8�$����7'%D����C �#�&wyce0��j[F��0p��#��� HJJ P�R��p%�V䋦ҕ7���#�Y	&�lG Z��qζ�+o�`PE�o��IM�`��&���`�,�>�9(�����"ɀ���Z�zg:0��`�]�ln;w��#2a���_��ZZ�0��	�ꒄb��/}�7�O�zwZ*6�L��׼�J%��"
���&��(��PxMOP�����. h�*Q��B:�LJH���m�U�".�csw/�_w���L"�L[��z�q��OFs`(,8fR;�%�vB�(L�� ,�R�t�����c$������4��Y�l��:e峬~KN��(,��LǍa\��3O'��F�p��������:����-*�����s�n@�V�n���t׆����Bc�ȴ;�J�����U{L�b���M?����.J��*�*�rc�c����]b�����ۏ��h|U^O�uPVȦ��$�-�4���n5��x���d�򔧻B@���x{�(��Mvg��(-j��K���x�,�ް������L�lb���&H~���`veJ��/�
?�N+��|O���7�(�c���F��`}e�JrR�r��.j�I{��V A;ZW��ҹ�J�.w��ͤ�����r�ً�w��$�����/� L�h;^E��{����?��-ω����fS�ym5�ـ󛻉,��*s�Hp�튻`�w�*��c\	��Lj�
u�L�˱�Q?4ï��"02�P#�KZ�����^D2�#�P�o��+s� ����+��P�Q	.���ҰU�-s�]����Z�S{�F�, L�A��7+�����n?t���/q�o׺X��"��V@��G���@�G�I��^z���yCBW����q�����}MqC�V��]xH3�FȊ��7���e%D�96ǐ�q;���:�i�ܫ��O�k�����~jzx��n�7e�.)ҥP5�PE��uCp�N������nEj�5���l��q���vK؀����� z���Qr�&jF�X�>�v��#�a4^�I��*sK[��Z'�Z�\����Wyj(F%�3�~ad,x̞A�d�؟�f�r������P!�g]�R �x~M
��6D*�����x���ɻ�a�J�p�VGhɗW#!�nR"� �K�4��Vx7�<��9K��6�%f�����V����I�\;��xI<K[����̪��R�����U�SAL�ms�
�,jm���?��|@�祍�/a��@b\b���x!%�W�h��Ds*���v߸�w~����c,	kt���̥Y\�����駋m�@_�fg�:;w�#�t����sI6j<�t���*VT�͜�>��.P��(�l��td=��2��l��Y~��a�E/���ʀF����o����x����X�q�u����'��¬�8�v[SP��MS"
���>
�˅�,����^�H�T|�1��h���) �|��7�>	��;j�>TJ��!�!�Г:��<<��.��>���E�NC,T��^[C�N�����B'+�+���
���yn�� %w�g�\������#��_��5w����O������a<�r���H�Ӆ`��^$�*-��i���)�A�쭬� HP��{�L�6e����L s�S+��� �;�3�$2��L�	|�e��4-� �	���d�nP����_��@I��#BK�0#v���5THӉ�yCnqz�x���0��e�����.v*��fI,my2°w��8�KS��I�ET��ɸ�R��Z��J�������Z�To�y!��f.�S昡2�G�!��f��������T�J����f�]��C̒�*F���z�$% �t |��H�D w#u�۸��^�K?��"n�56�"陛^���L�^q���j~!Ԣ4��3����? �R����S���槪����n��]���(����o{l)��r��,����{�G7M����LMA������{ap��^�R�!d����\�������|gfy	yw�Ҙ�Hb���oiX�*��?ϴ��H�&�aJƊ_�nM���_Ce��9�-�������L߻i ��M�X��C�q�A�A*��ī��$���w�^/��x�P@�����L[���L�@§D���RF���Y�84�F�(S�� ,`�)�Ӣ����R}���B����%2?XK�d'�(H���Q��U�d��o�����w��=Cn���m��0�q�O}�VCwϘpn�{��y��	��K3~�]�E6��Ё���vO�RB�4m�ف�aH]��y����3��FՔ=(�-�������#�=g�y����?���Q�i� r�:P�v����K���HwĉVd(V�̷��u��1o"Ƨ���J�W^ցᐺ��x�ӄVi�L�z߾����rh�ZBnAI��d �B�Bo�����{P0֨�ϕ�j���5Ϊf)����uY�	�-ݨ�,*+ػ�����!H�uk��!z��AP�'�<�ǂJ=���й�]ZX�G�A S�/�k��o��	DIp'a+&���
�W��f.��t�<~E,�?�4��|��`j����{��l8�K֢���`̋NCHp�<�T?��=-�7F6V�w���(Ĺ�u�ҨN>5$leZh�|���bK:hĦ���k�Z'	��l��'�v���K��9J$��OVv� �{c�J���8 �es���1u���k*��W	��D�{2���g��@�'��M\����O�0>_�����V��dk�nD�����M��`Mt�ݛ�h�p+Rw����S�adE�b@�dR�_F@M�܊��$�vZ�?֘G�D�Ѭ�:�֡L�D]���gͻ��<,c��^�8��^�6VU)���L�S3�om�u{hN�s������L��v�9�0lL�
��9�֨���lN���Gt���˅��A��NW��0�J�h f�
S����C����e/ ��KMɊ5
J�E�/�a���P�Q�e7�z�[zE세��TC:��e�<�-T`n6��U�����#���ݠ�$h�ʇ$o����#`Du'LNs�⿜`ot�=�k�#�ǹ�蟽02�&@�C�v��Ｌ�?���Z-���[�3����y>󋑹�Ә����vCЮZ(K�A��GM}ޛ����6�'����ƅ?�?9^�2&?1��KE�'���\���}|r�"3�������
�^�[%���ĺ�-�?�Au	�N$�3�ΏGuD
xY�d(���3���Ɏ B�y�9�N!����U�4n����ťu�Q��{Tp���84�*����N.�h-֕��t�IJ�����yk-ꯪ�����!�)�(�K+��秈3#��}�����C��g�n�l�f ^�HG�@8=.5eJ����P8�����g�z~HV�����AnF�;kA��� _P�]%��q�G3���=����O:k �gD�_���9���J-��7�����Sa&����E���$\T�M��,Ε���@?��lHYoO�p��nL3�f�$V�IO��p;�ڇ5�D�������&�Y]�b��#c�w��q�W�MO�!�}�6G�(��mn�9p'�EVi�>	v*��7�����^U�c���	5I�{��Jq��Hu)Wue%y�]�6����2�t,��iu$�<OVͯ�v"t�G���_�1>p�f���$P�r�����o�M+J�CX��|U��<¤o\�}�d�Q6�l�������j�dI# �*�?%��)'��ȝj��9u� � e,�ٺ���F�)50z��uT)�:��Xv"<A��և�Of�H9e�b�\w����������3�Y�Qt�����I���#���Q�(������ ��ڗjv�^�_Ur4�B�/ac{��*�5�COx��AS��>�Hzx%F�����GD+��"Œ��Į�I< 9��R��fN�䷑ZY����9���O��V�2�� 룥TjK|}��B�D?�
@L9Ih��v��{��X�k��t�W��nV�h �<�˔1T�q�׬>��}���Go[RJ�GtMB�)�C[�ak:nv����ܯ�(�x ����y�aɖD��I�֡�ՙ�Ʌ1�܅9F�s�S�7�����~E|4���7����Mp��
L�qff&~��~�8�����h����#�_-��@/%˝ؒ:Ui��N��.���c3��ic��G�qX+���x��;���M�I bЌ��I�#�^u⎗��s������X5�¿78+��z���-Ƽ\�V�w�=��Mv
NUjGG�oQ7�>���s��.]4V�l2o`�P��4+ӣ�Z�^x^������vko�����|F��
4:s'<�����Bs��Y�¶ExS�4��Lk���<$x9�~�Ԟb+��=�^�x�(�V�\�N$�������8@@ܨP�X4"q+\bY\n���-�0�S�C��5@v^�c�z���(nx;U�eY9�'ܟ���~��pK��z�	-��[��צ��`�՗>97���>��=��u	j������0+
.����R���M��FN��"�U/�y�|�߷���O������"��j�-��tҧ�/����NBֵ��79�O�t��"8u"Z�H;�� �w:�g�3ti��4�*��8�!t]���>��G����<k��L��y�k�m�l͌_�U��Vmj� �E
�\Ore@�$Oz����I���q�	~������V��`%�䢒��[<�,��ۼ%);N�&��t��[8�!H�vG�B)U����.�}�����ɶ�� �[�+8>ױ$�)��4lA��*ف�+F��2��~�K�,�N���|����)6t��eWA��%��P�~�gZ�w~��|Ħ)�Ҕ���/�(g�l��
�p��3�L޻9hMÐ��� �����0�!�1�6�:�Ț%gp9�Gw[�!Ď�]�넫B�C{F����yZ��B��u��g1͂�/���H�y�rʰf�\J����z�l��F��ߓw����~q�$.��>� #����Æ�3�>+��]��7��f1Ṏb�<ψ|�\w0`�Fڱ���Sw�>�G�	�M	��y��"s�o�T�#X(hY:q��)PF2�3�����#��0A��F��@eUehz|�o�Z�I��0Ʒ��I���ɾ�g��oy�������s�*m�� ��> � }艷�$���9|N�Q$;Id<_xW:x�ȍ4��"�3�����ؘŃ2�
��ƖZ2]=o#4S�W�ό��[4���2�y��y�QR�n���Bi��sk���<��;��'�s���J.$�u#4�B�A��znzh�f89��}���Cc�w���'�3�YDA.E��3/~�<� ���������k��d��-�qK/7�������\�I<1�V��k&��@E��òc!��B�I�`HϤJ$&P+o@��o�枕�<9՘z�Mg��o�?Ϲ8�r�!돓i��At�4R~BN�s��O�5����29(Dk(~����d��( &��C�V?��-��)�{ͳ��t��)�2�mtG�!��ך�-1,�iG���~� ���6�U`�t����I�%�0�r�.h���_���썗��P0H�<�KԶ��d-�L0S�B�N<`����W|����V���n�
2ǘ[2�F���� i����[�_
#���b�KG�&�~r�v:��^�~@Y[����-ּ�̵�R�A(�|�F�ř%V��R�n9�������^l�D������Z1���)�k�!I�m�}�i�*ՠU��q�®�������~��c��E��lEx<��᭄.�I"4a��wZ��G����5I�vv�%NW�G�x�����q����G��ԭ��o
��L/Z��-@T��1��/#�����k���v�37:�I�}q�Σ�a�#0u����q^�L�Lʏ/m�a���U z��yt^������a����W�)��񣰱���R��mY�W�&>yg��T�=J6E�1T�"����+@���v��,��������_ݮ�ͽ�Iy �[�(_=�@z-!<�O��+�>�f�ġ��E����]T�6R	����&�s=����!����[�,y5�_�)
��T���Ғy�U�r%*��x�V$1��o�3��ufX�� JAzj:�YrQTa�!DT����An�Njں�<o�M�[���GQ3���ЩSn@�,#�i�iاm�Z~&"�M��i��ϰw���*�����1�ꎯ�լ�W��'퓢�ޮ�	A�3��Oz�������yG��w��<�[�d~5��A)�u�4���l�
���ۅ��d7*��_�·���~hEڌ�PQ�����d��F��v��]��k��ҟ�.=��GQ���A�G"�����Ze�e\�	G��j��h�	:K��W�_b��1�|Qy��P��}�Wd
y�Ò&3W-:���;�,T����w^ ����%������%�[걟	P��m$������Mx�=8Z%����m�?a����o������+�f���'QP�>��-ALWK���!+W<�鎹#j�(z��=��vt>K!c�fm&W�N gm�ߋ�(ySZ�����ٴ�츺��۽p����OHӠ�L�=�g��M�-7�kϛ�&�m���es^*�4|��p�&�2&������C��������ZŐ�|g�"�t�iZ\p�k�x�tc�A��9Ӳ	?�(�+`7�I8W�6xV������p0*�*rۃ0�j�$����<�Z:z���,[��7U�4�0���Լŗ0ʪS�A�79Yd.c�%�_sw�Z����P��Zf@���Ȣ��d�X���Q���qb3�œ�k�d�E Vb9hw�݌����F�R��6Y�/b6��B}nfg1��f�N�ibnV<[�9t{cTRi(P��*@���q�|�i� �~^[�c�����SQ�t#�A>zg����*��1?k����8��W�aS��dBUtBʾ=��U�*��M�a��[ύ�zs�tf�A�RˋR��!�O��mJ��ν�di#�*����Dr�=�-��p��#��_1)��Yd��D(�|�xZa�|tʽ&Q�8p�R?̣��د r-U�Ƨ]$�GU��5�X���Ih)��3�L�nu���.�z���BfR�Ħ^p��R�::��F���%�&:K���jo�ti�Џ	���5������=6���𡹅y���Y@�i��!{�Rw�{9�����Y���Ȁ!�D~L6���^�:xj`���؀�w�-}��3&��/P�����(`(𴧰I�b�z���fV?E�l�YHM�CCo�Αx�u7�d*/~��-�@�r&I�
�<�"g�&Z:�@��F�Xi�d��5Sm����Ѩ�n�i��+x�MR^]�8�I��駖��d?�"�O�s%m�5�2��t� $��������+&0t0+3��dj8)&m1��9�3���q������r�>=D� ��hI�A�qV�#����b� ���=(�ږ2b�b-d����@MJɃ�.��>t˜0���s%	��?���ŗ�E<�zuM�)i�3;g	q�Y�X�Ѷ�i���'?5Nk�y���h�ϯ,:yY��6՚�w�s�$���_�>����b\�й������^k}~j���G�\,N���a�&�(� C|��w4�R�u��C��#� ⠩Q���[n�l/+�v�����:�;��{_Ծ>��M��.�.-��CQ��)��1x���}���a*�rR�#
V����E��/�hՇU�J��=�k^K�2�;�� ��m2<@3=R�=�R1Kư�:p#��)׼��Gd�=�!��i���`�B���ȵ��F������x!M�ܖE��w�߾����^��t*Q�I�	�B�EF���{V@��A61{����O���(ę���Y��8������ �]�:PT"̧F��bԀ\�������zV���b��(l�QQ`8K��<������
�N����e�,�M)�}:	�M�Q�N�{����}�n�l�����g�R�-7��g*��S%O��r]9ut�Z]��F��?s`�F�մS��
�t0"��`XD�%i�Ov��{���s�����
�께��b��;O�گ�+��>]Y.�/�7�e�����Х�>�ǌ�W�5�hq��
~ł2�/-Jc�@��,l��t�E@�Y9���A��Q����$f�N�l�46�͗�>U�}�1d!�prB7�ݤ;���h>�@J3�ٗ�-���#����<���<�+��T�Q���<yk���
hH��e'�1�u� ��lnhk)vmg�
a�b�cG��E {�b�P��&��(�"�ھ�� Tb8p�G���V� bSɿ�@ٰ�%Q,c�yk.�b���@
0ۺ�\�9큊�9=�����K!�	�7�,�B���f�W��u��|o�R�K��"���7\�+%�:�u�gy��\4�J��?�7ܫ��}�j��"i��<J�Ϗ,.;`WՆ���x�*�󲀣�];3����(�LpBHa[P��,���ۮ�����lU����[���\�'s��ig�Z!�/T.�?�u���V��_��C&�9�$>�w�<�����Q7"2 ���O8���s��x��NvA�*�z�Oωk��<$�?�sB�KR����U�H�K3'�AsΌ��@�|͓�q&\�l�`>Нɖ���\��	���,��9=]^��F&|^����..d7��G��� ����: G�ӪB:Ř|\q!��6Ҝ����K:��U����x�L��K�����Y�u-��)�F�#�bQ��u1N,�[�0遆!h$�.�b��Gi%��T;f��������{ʬ5����-ٛT4U=Oo�������� 
�߷h�+~?�֌Oy����*�n�\E���Ra���7ِ��v�dw��K��fu���.�v\Ӷ���"�����&�/�����������"�\�@��L�y��3�d��)���{Q6��(��M0t����e�D�E}O����)�b�ĝw�y��>�HI��ՂnkC�j���X�v\����D>I�{�Il���i�>���J���7S��g�@�)���@!.ݥ�p@:2=��g����6K�*��}ʃEb�'m��F�&��UE~�rb�����U�ל�X3���Dr�p�6N�5�-e�e���t�ќ�-J���y��3x4Q���`���=���H�.tG��|梈 �G�������=���1�'�6���"�[èjca�|���>/����c�*�ƹBE�Jx�)����d5�Ϯ����֙�V>8aX����th��p"-����]o�])JXFWb�?ߟ�B�W5�#��H����O�����;
����l)!��7����ՄF��f��$�\��f�A��ca��{���`���S'��[1)ֵ9񍣾��lk`Gb�l̏�bX�~����J�).��";zgtv;ROO��T`'� ���IJ����&�m�g?`�i����&C�W1fx���/��㵅;����͖��Ԙ(�|i��v���M��S��1���Z�~�=`
�4���ު�M����@t�K�r�㜢]U��v���XM����N(�Q���}��em���7���z	�|<R3,�o͂�ջZh�M-���1r���{���ژo�����p���P�����{+6����j�.��*L R`}�>���,æ�R�UnKz����Ü����R��p ����$l��0 q������e룋0u��{�>�����h�f��*[!��O�"!�.}���#1SV�0�q����lоӼ��EAj��K;ݽ>�Q���K��ci��r�C�Q�?�=�lb {>5�2��L�岇;�"���1t<ʈ䗾I�)�F����� z#+D��?��~P�8g'��¯��k�P�p�7�dx�&8�Y��4-�.�z�U'��)UĿ�6��5�;J�������Ʌ�&ONĭMJ�I��� �L�1�7���]Tc��������(�j�����D�4/l<	��[d�e��2�U��7�-SK�5�7d������:/��1P�zqˡ�s�B��]�@��̄��	���ŧ=��;��9�wnft䤗������u4t9�z�ry/��z�����]�����q��j3���ߢ���!��"�����J��Q�P*�r�5'�kH+m�E3���mތ�·��"Vgá��%�x��h�y�HN��j.^S��-)�_�۲�!�%\���#�C-$q�!�BI�>��b�8|�:u;:nO��$�2a�:�e���x���a5��j_!zG&f@�3������=	�"ϢRʊX+����,�����n�7�(s7�X0%��9B<�*�� ����.7e��� �p]u�ZB�"��ƪ�DiCY{�R�
�ɥ7YW��Ow��1�鿋�mp����{ZV��?�;�_�����JY�D��8�:ׇ�~g�\�$�r���[���6�sZF���5�_��(Z�������dEO�B�Բ3\jۥ��PO�I�`ExN$|���>�ސ^�a��Tn���3�L<]du������h�ʉ�����-�{�h�7/�!*�W�����N]��,��¬��� �@mp�Da��3�P�!&k�.��i�&��~L���|��
�,pA��W]T�-���>,>� �ɰ�uoS�v"<����;�y|�5	vBm�Ӝ�K�.v{�VyѺ`2<��@`ᢪ܈���-j�x6��;C��\;�}^����#Ӷ�[��¿�XWrOO`%	�󤔭Y�֜�9|<Ixw@jQ�-������
T����
