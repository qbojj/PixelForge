��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0F��A��+�D��_UOLy��H�{�i� �뀔q��qLU^�F����;g��£�!���Ç��F[v�G�5f��#�m��/�JC)$:zï�C���ƹ�xc�N:]o��Y���f��?�T��l��b�U2��h���Qy|�Ä�%]�]V��i�h�E��fm�ԣ~E)~kx�b�HX#"zw
��N&n��֯3 6S���5�_�Y?}v�����E�F��,��l�d���ӵ1�3N�p.�P@�=�jCO�����C�v��*w�N�(&�>��WLɡ�T��%V����e��%����z��U�$u
�QJ����0m��v��G����0�(蛨?� ����ӆb��4�.�g��1�}*m )o��?ˬ����y�@j��`��#����Gy��ش�-��%8 +y '⬙���mBn�u�R�Wp��_
���BZ�S�#7F��'Qy�~ʌ(��X4�as�l�]��E�B�hY�x+v��O'*�wϤ?��$���mU�����<�G=i?����aC�����PIψ�V���$�]�&F'[@������<DV�����y����N�2�|;w��9[t��7�0VQG �� _HC��"�}ΦyurN-��]>�Y��kxiQ��k����g~0�}�Y7J�8��l��e������{͈����k����Y���&��)`�:@1����[�;�͉ULJo�F��^�Bp�3��SP���J�z���d�o\Z��k��ig��/�=8�������R9}�N���p��2��B`�z;�b�JTC`�qg��l��^�""G@h��2`8����s݊�֜zQ���P�+����}7ޭ�&�,�͚QO�S>c���\(�>8x�c!��3������, ����/�����~m�C����lW����;��<g�����	�ܪ\���.8���J�k��yN��t��'����K�V�6�}�l�	�Ģ���^���=��-=�=�(����00@�o�-� #r&���l����a}�7�O3�D�mNq�ׅ� z����[]�Q��1X�3ϥ�X�>+ꮉ��'��ԲM���� �E�
�����xg������K��7=^��O�����4�t�� �����
�F�##NM���j�"������{�*�ݹH��\�X��� �7#r�:��n���Eg�������ҫ!����ؼx�6���vֿ��fb�1�I�M,L�d��ô3��XO	��
��%�l�,9h�M��xAҿ ��������.�3Ê^�N\���6)��3�VN��?�S�k�w|\���*e��p�R��կ�W|�fܠ�UD��kJ�[���3��,N������ti�~��B��?l��})
���+�s<3�F�
��R��ߋ��wW7
Vd\p������|���"0[Y;Ɖ)����髴��H��6�*降?��5@m��A�,��He5�G���)�L0F��� +Xi����Ex7 ҃�Uf^CDy��?�X�29����f� �֠IsOkN#�"a�o�m�;��zA�)�{�ߞ��Z�Zf$a�9�=!�J#`�yQ���	���r�C4�Op�R̈́,~!�j��P��Hn�u�X�Z]s���QY?��W����0��N����� X��Jt���k1Z���z�{��zq������*�Q�7~| $��:����:�^��7�Ǿ�|OKB��j�kzN��v��;}��Z�����;u���%���	���Ʒu)�Xu���>{����"�k@���{�������6���}���]�G����[����v퍆�#SKp~cn1�'~B�5�?�d��:������p�@�W�6���P��Eu�al��W�Z�����w���E�[�t[Coj��Ϗ���܌�)j/�C�%�5���=𤢑��@��Y_�M�*�s�k�w�5�8o�[T�n�[Kq\��#.jYJ,�Pd��1=�E�9���<)�<���6�����l���/+}'�$d�<�\�}�ʣ��N�
{�?�&���XJ����*94ǺIW�Ռ�g;^:�N��8������i���L��9��9V��^Xf-�/�P��om��ZyU�����Y���LǢͅ&k�f�~^�M�*�汽�'��^��q�/!���V��I�l�d�I��QѕYv��.�tvh��o|%Z�����I�9G��* �+ҽ�� �yD�$�&�Gr�s��tN���A�~�k�#8����d�Z{�+�a�-5L���ɦ������w����=�'bW(7�02�1�}��be������j'�At7%�י�G�X �ޜץL�XI��4*�ZC��x�d�o(�l�`ݔHV}	����8v��^�L�c{��bǑ�8ґL7��*�ל�x����R�[>�@ї*��^��l�{�����#,�V\�������:�K��kf�`��$�du�)��8׻�%G-H$Y��E'�-�o�Z7�`�2	.�o^t=�vf�5Z�y�`m��J����4���\�wpЄ+[�	���� �ؙ���ɧ%��8� 	E��jb	=�l���K�����\mX�����)�
C�B1fK�e\O�����|�Z�yv�$>�ݺ
�v�I�N��p����>ꔝ��~ESN��3�I�l���+5���]���1V���I[.RI���З��Z_��V����񖥯&5��kuh)�*~�6����S)�w�[�V���2]����%~���xQ�D�v=��1"�C�E� D}�����7��Fp���*��Q��xz�����|Qmj���L��uP�S��mt�o=@�X3�Qg��0<J˔��U����UO3>Zl� �h���+*��.�:�Hֱ>x	j Q@�5�V���^X�P�C��C�c�Oc�PLvO]��^�L�`�b+U�s�oڊf�@��G�'����V��Q����3�]i�wi�|�/I���rl|��S���8Fx~z��t��dڠMϜ���9�E�֦��P��SԤNr��1"X��V�T$ՙ���˾Pa�왩��(İx,����F��bw&��W���8ǽWݒ�WE���Z����㼾�ý~�$��&�9�lu*�5�"�5�3�m�z�Ю�֫��E��-|�-lF�X���0�.n)�QK�Z
~�W?m��bR.|��s0���:(���&!����6L�"�?�&D��Z�t��s�N�m��I%��D�m�����Ϻy#�y['���x4(��e�]9)x� ��-����D��h�e�_Z����؎c�RH�__V�L�hTvO�)�:�:�X;p��+NG˜�]�9�����-��̙ƯfO�	���1��zv�`�\��_(�j�|�mG��f=��<ZE~�T>E���4|[hZ�Q*�V瓛*���)�E\c�@���@��A5}�o�Ƕ21���H.M�*1�ܓI���_=�i��G�A��v4R=���:����Lg���O 9�K���綦��6��%#"�e&��B�l�0,�j�;���d�D�%�������;QUz9��A��Fz_	,�ڀ��c*f�2#�Z��?Qδ�^�+[k�5�
\]�晓����)�A1��5�=rl	Vd�0QQ`*r�/[�yF�Nm7��hJ''_��XA�Z�ߜ�BD@��^i*`ϯD���I�"�sM�܇c�n�nKI����y[8�#���ҽ,+�_W!�WӦ8������L�n�����X�=A���5!c"X����~4F6@)>�5���S�N�/�� V�}�������D Ժ�^�ql&��#��yn0�k�釒��O�>C��rgCCO!Yc0�T�s�|�}��1��V¹Q��w�(��S�a�+�W͐��u�ƶ�fnl�|z�{u 7�l�䦛VT�A�#�ؑX���Ǣ<� q��е%�}bŗd#�6\�o�s_��k�dJ�o�uũY�B�3���p�W�#�b�gG��ɿ�E;VÅaZ���P��ER��߀�аN|^h{�h�1�XdG�����_v���(�
��"'��J��5!�G���?z��)}.�����O2k�1�[���AeG�4鷟�`��=U	z�48�Zu��U��49��#Q"_���R��H�R��t>V:ǳ@���wwmR���ULZ1�o�'��Mwʰ���u!_���5x{��`�C��>p:5I��'�a����%�6�̙u������J�qcT��~v����nF	�*��AU���)P$[��O��?V�4�^��Dt����%oY�+���|AL ���X�~G�H]��$����A?�@>�=���7̒Ȏjo|o�t�T�C�����
��s�,���M�f�^�Û���{�z9ڵ���S^�a�n��<M�ſU���ܟ���Slnu��J&���	��}/��M�C_���̮�Ή�r�Cr!+���lBg%��W�aD鯴h!�N��`z�"�O�1ыWE��V}y;��Q���'>�ӼL�^%8�R|D}�&޷�'>)�ǘ���Q5�<C^�p�BU�2W��}M[���c��z�[C����lP�u�S
��P^s��K_t�t˹�q4Ic�X��RZ9�B1��C��^?����;k�ڋ�2��6�Sy��U̷���eɁ<,�}��0�n��[��'��;Y�T?�xA[�J� ��C���Ku�в?��
�`�ϯ�o�&����Z9�]��
�~���0G����L��Zul��,3�3Y�,1t�Q/vj�B*Yj��n7��L������1�uZ'h�aJ!6a.G/�o�4o�Mj������%���P�4����#����^V��D�a�3-�n����V��%��tܥ�F�E瓠�9ܥ��e�!�0�Jo��Q�������!���	�!�����EmZ�[����s�/}Pxf�MT��:F��b5GЯ2���o�)+*U�[lT�F�.��8��B�W��Ӈ�;�
�K<��$qwf�W���!��626������9:����c(�st�"��`,��@_���+R<I��M��������S���1��P���8l�IE�ұȫ�Z��R����PT�X�zז�1�ܘa�8��'��d덠�iv�������n�*�"<Q�����G[��>�T"�ӽ��gU�MQ+Q���r�dm� \��W��3����3��:(�F�U�e��a�Ƕ������l�<�d<1�I��뗣���Տ�s�w��I�JF�,SK�����!&�����(�#���MV�!��>匌;M�qy�?��A��ҵ����]i_
�-{��~�x����l��=(�WV��6�Pt�����ǔ셱 �ۇ�*�A�{����F2Zj��]��������hǄ�_x��6�����:S%>$��U_���8�u�1ζ F;a8����|G6�z%��~�b�R#���H�O��O�V0��G�� �!�F������nt�6������5�X���A�^nQ)�&�
!��0��A;�Z�Z0����n�1�[��d4����G�'��`iD|���|w?ן����W>�s��S�I�Ђ�cU���[B>RwrP��Ɓ-k"�bĭķ���$s&3�槑c��2{����iP6�������&s[�û`�7ԛBh���*�Lo^����ɤj���gvK����T�0D`�fF���^֝K���L�-x�sK|�K��Ƕ��m���t�,�4�8�;�bLת`2W<��J�f4<l��TlOzy�FS������­|�ݠK���[�c�����,~���){�݁��q�emW&��ȷ9}(ڻ'#��Ď�|	��S�4�\P��fl��g�m[�>�m��)NQP�GA��i���M�(d���k�ʘv\a��ER�a�ŝ>�i�c[�����t��k0�3lz��r晕�QZR�I��ח��㩻�D��L�����������	)�����B�򉧮�2�IV4�gI)��A��v��F�5���8�AyM����Z�:�Ez�=k��e	�Q��?�ꎉ'?��~�%��(��$X|��ք�fN�b�=#�Z�z�M�A�-L�{����<�g��(�,��Ty�a��0w�	��
wGZ#F!4㱼���Av[�"E�F�>%#��d}��2vEU�G�	��5t�m��)�7�>D C�U=Pm��Y�'��s�`��r<W�ц=ϰ��⁘�0#�C}�`<��4p�-���e����tx��»;�_����[��@m#�E��R ���96S�����3��j��?aV{j�&_�(q�3�8l�l4>�[�P�Xm�ⲭK��C�g��a�;V���s�<I�aOm3yq�k�H����Ux}$>���-"� �<p`�����/D�+� O���蠺���ћ�s�4/==�+u�$���|�����ntq�8H��;ь�wdy!�{Z��d~�I�%QG�\s�̦M�e]�W��Z���!`'�A��
\��>9���ʃ�ǁI���ٛ��5~M�c滇³�}�TI��ATl5�%7���c���ș�a����Tw�)9��V��NY��n�Z��0ة9@��g�	#c'�1ڕ8�[�a2ܓ�A��N=<���"le2d�N�JgM��q={+�s۾T�%|�@�F�:��-n툹�G,��sL��xX��B�rP%z#��o�u�p	����)����З��[./��ɑs����}/J9̼E���{G�A�<�$�e�-�y�H�^=tNiN�w����\���[���c-#�y�}"���KPF;b!x���k,�Na�B��~�&C��q����f�s��r��2J��_���&��=�X�6��r���]��Tըb���Zm�`z��Z��?]*��6M���gڒԭ��8��|C�|)�W�)ݟ:�?���v�z�G]�?��~4j���X�V�<���v� ��jtx1e�����ъd��ҽ�&e5Q<h�P����d^.�-B�ɷ�j�K��c���SV�U���w���AC��)��輈�gO��*��	f<���\N���r�jH���k/1���P~)Ln_L��ovl�.xc&mYmL�b��1kPE|��,�N �j3��;��%�I�mHG<��t��<f#��ϩq�����Ƶ��(��@�g�y��F�č��\*�;/��6�/���5�>V�g��{�����R|&�+S+z)b��	4.g���զ��V�ؽm�gs���Bݸ|Rt�,�Z�=*Uf{.d7N5ȉl�FO��(�j��0������q��1�>����c��Tt~�	>���-{.����D}��}f����8�؉z [��xA�F�b�@�r
�Jƅ���[��׸��4O���������6�8�'Gu�~�F�9�នG���tS0�Ta|,ۑNF�:��v{$���
��3(eG1Y4�b~�=0�6���R�x2����U�hU��2��O7���O:0�9s+���̧R/Z�Trٵ/߈�2�����Rq�_�@�S]�JEL�zxK� b���!w< E	�����7���5��M2����ZEU<�%-�+fB���x��c�� z�j���i���z?���W�6��CT���o;�G���09���K�nV��I����!qK.�8��*��~�m��p�*��+����|�b�K�@�S���(e��r	EI*m%c�`P@ݪ����H��5n��@�},P������E��Z]���p��d�5~�ۇL�ā9eD�tT-�4��"ηC��t���Sͮ��[��k<NC<g뿗�4�T$%B��d A.���x�z]��^an���믎t�����&�S�MsM�0���p�R����i ��� ��KJ>���ҵQ!��p)��@\l66�qz�Y���eLe�#{�%�ag�o��څ&�`j
�/Ҥ�TDq�ʵX��iZԂ�Zt������寍 +ԩ�5�VΟ��D�֠+;u�s�	d#����'Ma	m�R��<S��kr�3ߞ��A�=�_����F��:4���~Y��M�V"��@4��vH����
�ˌ�ЗDқ	>�E��GI���o~��J9Ys�32��� �#s�^�&O�
�������~\�_��*A!V���l�_��9qV�)�!,�F/J�48�!="�0�ծҮ`X��;.�AY8��2��G���:�K��j�.�˗�=1�����~ØXg��RN�G��3�Jin�DV���;�e�U(Or�2�D�ȭ�}*s:����<<;`Bӆ�P뙥Y,+9��ƙ���?cC|>�:]�;x1�궉?lNB�A����(�c��B0�Uù48�Z���'=IT�/<�b}�^�U=���O�2
�|���g��g*�QP�?�������jcH��{ш�Ъ�v�+���������
��?����q��W��I��R���	�
#8,�<�&�	��X?�!��m.!2��n ���6��Tx�V̩����g���_�ҙz*?(
oC}����D�"��6ioޣ)	d��HK���|R[��&��`�#���2.=	�K:s��g��ٗ�(k��6��"3�!$�7iX��M[�	�
����(�M�L����u.���R*P7a86r�-ۢ}��w��l����H���K~�F�^!�����5Sf����0
��B��D�ei?�#�2�Q.�C��@Zl�f>ul�T5�`YN��z��^����a�+�x"�w��]��qUQ��Ȗ��K�3��MN�j��v�6~k�e����	����状���ԩ�R\��k�����η$L���)%��ħ|E7uw�㽚�|O	:�.&:f�Pԅg����}��T]��2ـ.	�t+[�e[FF�(	�x��)=�E��O0��a�޵HsZ�)f-�u� ��'��*a� �~5P3SDOe����h��� M!G �↋2P�6'���+u�ϱ9�\$1��=b2o'1D謰ع���lzf2�7��& c8�j�$��
و���H�-��ڙ�ќE�� ��M����:է��G���� -+�o�u8ȃI��t���H=hP����.ҹ��jB��-	��a-酁a0 �f��l7�v�,h(1���j#�ϪB�/���p�����6�OS��K�y�/���5��JW#�^_�D�e7�M�J��{�3��^��gl`�?Դ'>v�v��7�J�RK��9y�;���j7�>�'u /,2!��|�XVw�n�Y�W��n4¤&K!��7��C]��W�HڍnIs�H�,�!-i�3"�а@7m]�����n�����:�1H�nj����H��|b�4#1 `�lm#Dr�/��#�� ߭N/qE$y�/�ԋ��䣍H$���W���j�sa�f�زe5]���A\�uOU��;�4������4�pv�<�7�f�I�b�s��"b�� ����u�A2�+�.+�p�D_O��� �ŒQU��Q9w�EP���������*� ^b0������7�_w�)�6.�޾N�8�^7�6R�G���x���w=�\��l����(6�������?�E�۪���(�zR���NԄUd=\�l��5��g�Alc�Kg�ḡLh
 �j�mzӉ�'��,"�m�x�d���E�&�-�V��F�(�_��Q0�p�3kɫ;AE���]��	�+�szwW�X����"�H��9�R��m�ej��i솜�dT���G`�,��-ǯ�#ȩY�N0�zu}� �\��>��3���]vi��T�SӐ�M���7����4լMʢ*2���p��}�G3g����]+�0�Z��H�@�P�s��X_�i�+��)�A;�K���z_�m^xAΚ/��Y�.:L�5з$zJ�� ��H_��Юn8�1@vD���>�`<�9�[a���Ԇ��t�T�4��b�p���k�mZ�����e-�i��:�
�mQw3ȜmR���X�D:�}z�_��ݞ�����f�h�!���޽l�Q�ڮ>�a��#g��\�qN�!�E��aLW�zz���e��baD!N�ϫ>���ʵ���*?e���ǅH�z���0�mu��cWKhRO�����h�o(�昅 =?P�2��=W��d}�BX9�/�Λ�TD>���<�V&�<[�{7Op��>8V��hN�v�N�wC�X�{���~�e�Kf��sq��c�"�҇�/~��Z�J��9����~$�Ѝ1��t>�e�;�b�"}D��m�ڻob.	��ɯыP/o
�/�Ҁ��B�
[�����[�O�t�M��5� %�����$��Z���r�q��cH��M|W]�0���"�wc������0˴�1Q�s%f,�O��GN0\�?q��aU�nvK�Fx�3�R��+duq6�҅��3�-#�'�|Nn�(�L�;7�sbn,d�h����ʓ��P�������� �� Wv�Er��n����!��:a)A3;"
���Hu�g�8�Ӡ7���6�����Z��$�oR� �e����-��{|��Z&	���3��j�H�q-�l����#!k �ݭT��Y5q_SS�nl7ϕi끔��t�jdRb��O�'��ܤ���s�.��X¼��|)P�Ұ��I�� ���_�\*a:)�N	3�����R�'���L.�&}&(�%��5\}�=�LH�%�s9/��z��O�X��ר���秵�,� 	�eu�{i�r�5ru�%E���+�����|	+~�H}(h�=)�c�Ȼʽ��!�t'Ƭ�n�ztJ=�/!��N�im�@(D3���p#��ş�a�o���K}�)RPBT�W�򎚎�M��?�g�r���
95,�h�� �d}� ��z�;�e	����Z�hmsn�v`Ms�p��o���>�wc���C5�t�[]M��>�0:�Q�����$Yj�� ��2�E������Q
��a���SB���h��#x�!��S�D�����Q �l?H_���$Nk:��gvjr�9��*�|"�>QE���UYL����B��� HE8[�������J��'�0J��t���Af4?7Hy�7�6�$���U*�0�܋��5}=�\�{Tw��������'�k�b�R��fҭ(s�G)/�ĵ=_Qi�-�j3X�\�A�zmI{���6�����[�v�0s5����G1&DK�X�He��0�o�����~?�l[s�I���y�D���A��$9���f�x���{�z�=NF0;glBJ�����C��;!怦Z�mC��T��ci9;t�����a�E5 I��@�<b��EN���~���ڒ��BC���@���j�
i���Ӹ?nQ����	�9���6�ͩ�H���q�5�OZ���r�z�AYBc4�9;����v���fqKsbf�Ɖ�m�"쨉r�p*iX(�.Y}N菱�yBV%�E���_�ͨ�4ѯ���4�X��x�g:���:��O�rK"S���1*>�uR��[?�B}��+�ӌ�lr���R=|�]֚�y�>O�Ӱ�5/!t��u����˩��ң��v�u�G;_z���A��������F��3[��������!$M���*�c���g��g�;�z�/{^��Z�fuI'��U܅R��Z�^a����բi(�n�A�U�͉�b_B��r�1��r<Ñ�Л��a-J��z��k����ף��g��8��:����?��zj�$M���!�G}I
B�>I���D�qD�c��m� z�>?ǧפ�в��xH�K��#�.�^Ek8B*�2��U�l*��3}�krU��z��Uq!����Wו�3Fj�!�������X�����\3�X�9h��}�a�D{8D�/�{�,����t$E�I3����iSf"LK2ś�E1t��X��	;�,fl�v������c�|	��
T}�Uޣ�G���|Z���0��L�o����QX�����WŽ�0D	I��z��46<��� dl��y%�_�� L�F�U";J`����t�� �U eNzg�v���^�Yq7\0�F�����+ú2�@�����,D�SLҋG�|���/�=|.��u!V�����L�l2R ��9�������}�YG�$c4g �o8�'ބ�Ч������]O-����(�G�gW�"��ŘV��i=���*�4��lqE�O����i��E�#"��F����WE�0�(��L�ګ�V�����fX+G_Rʙn�3kR.�a���ˁ���d��������MB)dQ]�7JV9�3��������]4;�i4
qW�I~� �kp:�u��K��r�(-2�8�L�~����:,D�8���#�g�x��byښ�x��A)��
V�aI���em����~���]>�l��lVF[&�K�EE����<f���ο�
����sJ��V{D��wF���xn'k�Bb�٩B�盼z��t�]\�u�'to�N��sR�s�@�kH=	��P�%ǃm�K֢�=Rx㦪���D�m^[�D:`kUv�Nf�'?O��O�e����(�k*X� B�D��\�#O:l��!l��Vz\��u}���i�����
��
��m��wsQ&`ɿ�D�f�Rm��m�9u$�,[���yy[��w���~����ێ=��Ja��Y��<����nޝ�T���V�L=B4�{�n8|~�����B0�I���%�$��)�ӈ�B?3B��(���a{l�f�U��W��'��;��7b�ns?}Y;�,銘����D!_�q�ᣨ�'��b�����?İ��9U�h���tX��]L��@E�Q)*",��?H����^�.(}a۝+��K\}�Ё��[�:j��lHZ�����Ț���Z��"�����-@�D�{Pd����Oށ6��*�z@|v��(iЏ�th���-ӉoHV��P, �
��`������ޣ[�l{���!��~��
Fe!d��m��/"l��`�m6�N��U���N3�1OV���Qw�
Ue���mk,����^�q�T\����j�B,�{�2�=љ�S<�|�A�3ro��3LҺ���m��P7|�$K���`��I�τ�q����O�Y��=��0��	��_����u�ԇO'P)�-1�,�t�
���H�S��-���{	d�T�����5sh���$*�{�F���ґ����q��e�>5�{hizR��p?���9_Vll���|�ٙ�I����o}�Ҥ�ZT`j��@�}�T֗bZ|UH��̭���_����s��N{߈���[B���g��f-y֑yQjQ��e�.���hC����� �f��ʥ��S<�LU��.�\O�ף�ú��3��#S�D�H��I��3.����AmkԂ�C�h�L��qF���:YD��($>5��`S��~n�ß]��Ѯ2��C�ػ\2Α gӡ��-qp�p���(O�ǉ\��C��9<Q�v�T���,����:�'e��1�꽫�f�����RX��[x� <J�2J
������}ºD���]��ȼ0U��r�)�6�̀����<�"�ȗ�u'E���OZz�R�tP���Z�e�ʦp�JC!T���C��l�[�U�V�����������9��\�	�!��B+�E�U�n]�P#���
��`</�ә��Y�wׇ7Bx�"���`F�h�Y�<P1��8�9�r&�W�;��jj�����c��	�G�c����nd"���}Z�ip|�"SQ��U��XT�[FLuX{M�Zw�����s�?d�A��W��7�z���2!3��d�� R\��U��¦�ܕ�փ�qb ���6SaD0}�!��1DV�!�{G�
�p �&�LJ��Չ:�$�_N�W+������ե,�g{�w	|d>��q;9�� �%���^�h�4�<��WD ���t��]Z���5���o"���u�dv�����O�� ��^8���bf��nl*�X��wj�����D�1L��:5a�h��o@怿��~鳁a|����(i[�
��ʐ�-��:%�y�t��*_�N��A2M���<Z�[(��!�T6�|t	5/ײ$�C��Pph�rm^	�o%0�	6*O��34�Z��Qi�r�Hw�:"�����֪E�0[[�-�����NR���u	�z7XïD�k�Sm���/v�(ǐ�٦OT=ҌM]��i��9_^P8 -����rxI���9^v4��րb*���^vdNx:��*�VѴ�lXy���Wm��C<\gg7R�`��ī�*$�?� C�`Lw��J��j���w3[OO7xx5I�~������kw^ޠ7
Y������$���ߨ���sn��A�p��۬�i&�&+�>e��:���H� �@��	���氢�����b��0��m����M�u5O�D�:������� -f(L��!L_�~B�A>j!��n�-������"xW�o��$������s�����oI���a����70�U���,����ع>E��b��6�E�y��'�.AW�qN���# h�i����<�)ݲ��&��34�mH̹���k���ǼV�4ҍO8�rI�Q����Ȧ��0��D+��m�W���pc9B�o�uO�6q�X���vec���cGΥH�?��:��9áґ�����[r}AK+��9E�n�p3���9�V���+��NMш�1��ځ��f��u�Q�ܘ�=&tI��%��;1=��x]D%�R�~���`1�i��0.��d�≤��C|���# 9�}�+_��ySLפ�'��p�x��w���fs؎.�l�H'��,H�>\;��?W�:��)�w]A���x[����d��7p�R�oE�N�T�,�H��N�o ���E�Gα�#���l�Q�������kAEl�y��v��7z�I�d�����ݠ�U҃��~ob�1bv��*%hi� ��uǐ��f��9J� o��Jz�Ձἶ
_(+��hi�����W=;9�4Mj~`ߊ�,���AL�U�VX���/w/��D�MZق4��M4U^�z�	��@oU�(���X�77[O�{���E�9P�ᴲD�z6��o����6ٟ��L����
�Eg���?|돲���-hX�bR�8=���{�vD]�iA�w�9� |p�*��]�n��l�P)�_ٛEu�=��.�P���w���M���8W�&��@|Q��Mmz��MX`�!�Q紮4������8E>�X�i�.��l!�rZ�D	������EM@<�8�5˻sSF4z��'\3��?EPݲ8��
�f�``�ܣi]�=�4>�)���<���Hw�h
�)�&�R�.�)H Rא?�p�!�RF[���2fF�7�˒�w�]�D���Y^��6���ӮQ�G,RyqA��v�pL*0Ӑ\ޞD~�ihY�S2Q+_��8�gqc�.x��]��Է�{�����E�=��q�Ƞ����*�o�������?�%P���_����G�o� ��Oh+[��(
�v�yzY��B����#�'�8k�#22J ��eL'[�F�ޜ��$�]��w\� :��E1w�)v�WH��Ʒ;'�k���S���'��hϟ��AEtzֿ�>ff;�����Z����	DG����N�a�}
�{�:�a��wn� k;���	�^3���*GF�������������iSʫ ���V��k��������6���*ڌr%ߏ;�A�
q�/k:����Aj�{�bX����|��+�^���7A/K�ŨBƿ�ؕq���{�Ԯ&�b�V�ÔQHVJ�+3	��x�"�~�T���cSe�F���.�U(��+���.T#S�	,��t�$�3��pPE�3(����z�ڬ�]�<�jG�kU�
�p��V��)�*�M+��1�xc�8�M�z���J}Y���M��(�Y��o!,���b��N`��/���<W���NH����<龞�9��j`�j�Z�=����^��&�|e�?J��V��=�����i�n���)0�5Κ���O'��/i�g��q��e�^���%�$Q��+ JL�m
��q��-��J�K��P������HD�����K+�]�6��ܫyB��+4&�W,Tq:���F8.�2�^`��P�Ml ���[�l3�����B���6?{��Ə�ѝ�*B.դ-Be0H��v)�����.�.W��S�=����O-����pN*�i�s���Z5��1��p��z���C3&h@]>l)�_���E5x�O�I+��`���b���;���&�ms�#�·	fw�<F�+9��W�2mIħ���5g�ss�jo?N49�U�@�ԯ�ԋv&�(��oE �L��h6�^�Hc������A��w���h�:��.��u�hQm�nG}�^�|��7=i�!uD�ґҐ���*�0��r EUt�d1��L�U��Ο��V�[!p/��Z�4O��ꔩv9"�P���m��M�3���0���	R��uV�v*�i=�n��	�ŏ��4�|~�X�p�F�/ 1�?�_����XQj-��M�Q&���BCu��~w�����Y� ���3�4��N�_��/�R�Ծy�)�08%#�x$�d����v݈��Rw�R�l��K<�����'��dt&r�i��%XD i�ŝ[�M����"ԛ]\��?�('��AHh`,��ur:�󊖸x:�z�A�T�}PmX�ar���� V�E� J�x�IA���{�킬�B-X�6n~��mF�h���`�?g��\���&��n���0=�������8j�(�~ �Ҥ��/[�0I5g�Xw���4�����U��m�(-ҕZ�!fڔ�y�澟�����Z��cP�$κ��g��٧��~%/�$�P, ��`:ɉ|����r"|t�+�X��ζG�c%^�勛��jj�Jx�����RY��j��g��S��'�*�c1���"�@��!&�V���!٬M^Ω�u�"T�Fb3Цx�!� Q��an��9_L�	�Z��k�,[�{^P!����~��lbClԀ�w�T�es���)��t.���ʫf���>WJy/X�hMQ�w��m;��\�n���.ΞȂ���"&{��c8g+����q��m��l��V��%��y�h#m*��tZ_�t\4{����bC����	,4[��&��������a�~��f�秨U7���\�n�*=��7��q<H>X�ڝ@hCx�W��(ԑ����(Y� �#3�i��]�}j{�?d4������u*\�Q� �6�~gm���k�`[l��V�B3�t*�	Zp���.Π��U���9�t�.X���*G]R1}��F�&�'1[����'��Y�)ԃn�:Nz�g����-��.��-�屃�+n��:��x�+�=����ܔz�C*P�W��`�KL�=J��7�im�S>lu�ωY���Ϟ/��r��x�K���ʅ!.=��<�X"P^��jFU(Vԧ�E��70��dЎ���ލ����PT���),�$��d̃��*C׆@�?�vY�*�Q�	h�g:rzg]�1;�J 5մv��9�<���e��1�8o�^4���G���z��A��Lc�RU�ic��v�c]Td^|�De9&�h=�Ǥ��Q���5F6B�2��՗��Ko�7A�Q�&� w�0O*|�qU^����h��w~�c]���U��vA\IPZI�u�e����	>o���|N~�Wf�G�O��Nu���/wD̈́�$6��^0m�(E{0&8g���_�]ؕ�����6� y�r��
����P|[z���r�ߘK	@�L��3�d�\N��8�j�tx�sӜ�QO��:��jH��:.;<-�Y��̕����\��y���
���8�m,����_[�q�3��~$4������� �jM��*��5�����x	Qxx��E�� �\).Qn��	��󼦧�Ocj���Y�zJ4��8�p�B�A��%萇Y	{������ϛ_���I��s���!i^�4�ByI��>'�����Z�r����0J�2Eݰ�	eE)���nد�=��K��mn�)���K��~�͖ s��{S�^�u���d��g��+^M��d�7`��~ap��Ŷ*��]y'\�6׃�~�Smw��V!�4�{g\o�G������A`���[�$9��s��%,��Gu�S�o��*�(W�3@+�T��g<�Z�w{��m�NW�j�؈�	���Y$�G�ڃ��y�:d��=�YKc�G+�෯l���ދyO�w.���*�ޟ�f����� �|��&�(^\�N�b.NT�@Su�Zb�z|
I�X$��ڨ�cJ�>�� Vt�O�'hUC���́59GϿ>�%�UP@Ձ�ֈ��J�V
�� ��P���j3M4J�*9�i������P��%y�Q��Y��~1���n�e&��,%+��夔�:�ǂI�����s���j�i:�<X��3b��)��79���_M��`��>c�8XA��M���`�"�y�tM���L�����Uܹ���#L��xx��;�фx�뼛IBSO3��a�%͢أ}Ϝ�]P��w��5*�A��.)������(�D��3�P^��Ý���@&��?1t��~Ne�*�� �m�*Xف[�D.�ƽ��hctr��S6�	M�=Z�N�0	�4&s��N�}zM#�BGK��~�Tl���-|�g
�
�@_�9Iu��jH,�v���7R̄ɳ3�XMEE��_0�F�"�O�~ٴ�3X����b$ �|Z �𵎢Cn�Ћ;�W�>�!d��I�aߌ	�Տ�".j�ө)�Fs��	������+�&&<=O1i���t�&�y�v�g��3)1�V8C9���x�P{\��0b~z��g�o��:J��I򤃬r��a�]p�E�ϲ���D��JCK2�RG��'������������vVTW?��tr477��>F[so��6����u5�8}���c�0.������hAn?R5C�kEm,#�mLN��pF���VV��
eeXm�R�u�͇��#DV)��C+ ��$��o"t�����Y�qD ��$l0,=j������C�<�*H��)�k@c��W�	 �D ǌ4)$!:K�����]l��#�]Tfo]��:��:�DB��8�o����Sp���!Aَ��5���$�J��#E ���	���3@�}������`$n"�RP��=S3P�p:�ed"���� X����j\r�# ��&��ܤ.�yQ}��'��x��K��\"ᒳ}O_��'�ܽ�l6G�~e��ؚ��+��T0׀�Xb�iD%���XÈ��ixY�gNr[�q��LCԛ� b�6���c0q֞�ͳ��w�B�Ֆ�Ԥ�c�祏1	XM���9UN�P���GR�	_��)����s�Y:�Iy�r �,��b��$�S3o*����
z_��4>��P�	�� 3�8"�c/ �*;�/�2�ʬ���=f*T;�����H�Q��?
��]�O��Bg���=.�Ƹ_'�$s+��T���K=� _}[!DeC�I-pr[��"J �Gc��,����,=���쒓"�r���I������G���㒯���A0�J�;�%�x���κ����dx�$D�7ʒ)�N�_����fO�y6��8�Y鍠�2�L��=��)���2��Rm��	�u���H!l��Xu�~u�ZǷ�� 9��;�
_�e[�&ʎ�2�̝����^^�Z@��3}�H+��6���x����Rj\���urzhO@��f����,ٝ��lX�*9TG}�Cj�(#��G3�9��B���%�Z��b�Z�<�p֦r�����J5\'<
�]5��vVB8G�Y��RM�I��+��NF�y�A@��/�h��1=��8�=`Aٓ�ɡ��mk�L�"/=�t�9�����;$�t4\�RB�W�I��Y.��J8��Pb�,t�Ԓ^�6J�}l���\ʘ�}U���÷K�j�P��]$� �0��[�v�/������%Y����A���Ն�2����P���:�ݶ�Ͼ��\7�kC�����Ou��ԏ )a6�`���m�&.�G�9B�Y��o� V}��G��J5n��ݽ�:g�3?�I˰3~w~�5�D�$B����R�	S��.Մ���� N��C��4��u�����S�@��U&��4��s�.GZ�\U#�|8�-��քn���#�@�o�
;�����pzU��,0w3���h�ג�NQ�U���AK�x�P�7�9����8�t�A071E	�C�#��Bo´����s9���*6�%�ٚ����Z��c/�sΩʂ��,��<#�%��D��e� mo����n/�I1��.VSUMXC�V�g��r�i~�Q�1�v�k쒼i��uG@'tӳ�Z��{� R�񲣫�7]���-�?5z7��+*�.#Ưa�N���.�Fأs��V �A�����(����R��S�;�Qb;ď�_9�?/�O��`�;a�x��{�`.6�nS^�ޱ��KOd�\]x��W��va���Ο��l�Cg����V ��W�F��6���K�f_%�0^�@(�Z�M遶[��A׏0^�
�bduغ��X���Ho�r �ogH
��#�k#2*l������,���9�4C�E�V�*a>���u.@��p;�NC��Z�g�J�	��X���
[�,���X��bfsaw��m�`��Bv�&����JtAzA���q'(�ꐇ�O@W��E�u���ָ�u�R0�G�Rˑ+��G_�L�Hd��*qy�E?��U�V�ee�I�mDo�&D*/y�0B�N�/<�L�M%<�0t�_����t�Hƥ2w�/91������z?�j�̷�>T�"�ך�0J�䢂RKF�WE�Bp��K�I��gьge15�-HO���g���._J��g{rG�Uq�����C4c4ڪ��^zЩ���9��8�s���'���	�ʹ+h@� &�G3�09�V�9c�iR8�B���f�V�Z8e�p<�&���i�;�G`��D��MW���0Cю/�������h�Wu��3��uɹ���l!�N��i
k ���*s��%�Q���,����@yb?��-���9 �p�=tLk65��@�$ |��,� q�vS|�E��/�v�Mï����o�n[���_>���O�.�Q#@�q?�5���Y�o��V$�.�Jb��R1B��/M!"��>�_��`��]y�ʋ��}�N7���l��(�ƚ�2�#�lѫp��Dv8�0�YV`���@R����o��7���L�C��Dye�c����1���;�p���Ӈ��S � �����\i��E�e�t4b%��7F��0���7$�͌�\���������i�c6��eL?x��ǚ� �T���	6""G�#�zreI�D�8�� �.�>��lVM!��	������c��W�����|�jCt���+�F��� �/0^���N�
t�w��.B���z�F�':�x�C7C�,u5~�^R�9S]�Q(�$F6��jUKW�o<Ղq��{����J˂���1r�wᇤҥ���l��!�Z�o^]d- O�[p:���W�M+�����S���tʃ6=��08�[N�_^L��qq��@������U�Sd��u�	 �4A��b�(��g�!�KH���W
,�e�L*x0zv�
�+hG���Y��Zzd�rl��T��w�9�V���͕�kۙ:��*�?"In�H����
�r�s6�D)�4��)��u�w\N���ߛ`x����M�5�-Yr��� �zZ�<��n��f
�QF�`��?=�B�b���0����4'lGS����`��>&:�щ�]Z~MER� ^��3�},3�bІcW������z���Tj�r��G%�eCQRMˎ�!])Uk"
v�#Ӈ�Fɚ�J�[w�� �W�WO�xg	�fH���xd*������㠂U�e����^��U7�g	�{L�3a8f�	G�o!� wc��A�����zf�u���)٢�ժcgr��O��"�Ikl�(����C��8�굿빅�?�Q�$��RW���ǵJ�`����q��/~�����6	�u��s{��&��5X`H_�ؚ���&���s�R��z&k�H?~b�E,cv֨\��W�C���GO�>�VP�z+������-�<_�q��i�Q��)�ƈX^{����""�;~�Fwl��@B���PP��Ϸ_r�%܋��=�S:��>]. ������*α�O�e@Ih�/T򫹛�DR��.ŋoN3k�q(�n����v���ж���l������Q�˂�����`�$:m�v�zgiB���Z��i�K��m�jF�Ls&�-��Qwv����t�<�yp�̷��$�A���4�$�[�U�%b���^K<�2��dKw���v�Cγ�b�iH��a��f,�}��#���9��gt����([v
Sd���)�l]ǈ�l�O��=B�Ϲ�d4�"�39��p2,?�`�?���Ű��Ŝ�J�D/�vH�
���k�e�/_ď��0cՅRq�hP���7�+�� >�s�]�4-BV��a��,�P��*7��g��w슅��0�C�NԊ�r��|��s@���n�3�?"/a���s�g���<��ku��-����~��x�LUĂ6wͻ,�oX�%!��y�: �D�8����a�q_ 6�Yy ����;&>4~Wݘ
'��%�t(����`�N4����7���2�;�9V������[O䥩�t���g�R!��>k���׺��G+�`G�O����4��-�w�O�Î��KO�?�uC���6K�h�\}�����y�Po]�oL+5�3a͎q305)$��N}�~i"��{��L�%D��R��eY�sRL:ʐ/=s�D��D�����vP喜�e=��1a�w$���EhlD���oi��Pi�v��hA=�I�W'�4��A�	��f�e�HG�Rj�Xb���΄r�(�`�rd��)��VJ��:[]�R�>�����p��\ӗ �ɭ�A-����pvœЪ��]%��nQ��Կ������(���Z��^Mκ�-���:�l�4��k��%V�^e9%�ذ��7���9�n��sQ�m�Tj��Y����Fb�"��M`H����l2�O6���t4޷�����8%k��Bژ��^t,�f�%I!�}���[p0�W�!�Qp׌�;��װj0���,�\*usFh�y��I�����ybVG�vu�m)I�L��\�m���΍�XP��o���'�Y�	"b����T��k%r!q����=˲�Ư �t�7�$:�qh�3��(^��m�>>�H� ÑJq�Ӱ�$ɷH�T+iq�F�J���_M�.��$�6N�|A��H�FsT����n����w�%�g�rZ9S}�����z���Ow
B �xKg�� .;����o����=_�s���J^p�)�lDkR�[�8��Uڼ<h:�R����
��v֥�����"�Eo8�f_㽠Ue���Zz�yȗ^���Y�����Ն��\����uJ�6t��j���;������� ��8��=�o$�������y[>{g�@��@��J�[h�!!��0����t㗫G����+�O���'o��Oz X�r���j$ ��G��$�X�2���J{�aﱟq��J:���ߐ&��c@\����?�;����K����)��*�x�lT�y���9�W	R��\���i'
���H�����L�3��f�5�G+֖��]��p��D�
 ��R�EG��02�î���?�-����x�vozU+���;{c,N�V��$��Q��H�`c��?�U�<̲m{���b����l|�GY��u!���'3�֗��5��X����<���2ę��}6�g��#�Y/�O�/��E��6Ԭ��^qG@�j�f+�𛪍?�v���>�#���z���k��c�����Nw�-�2#�`���	9�(:�W�%<�*�_Єs"yWb~�W~}��YQ��#�v˳=$dYn�ږ�"?��j�ȠF_���.�v%���T�@W�ne��0Y̨w
S� ��춞}�y���u�G�>��؜s�;Y�iٌs�n�YVc��MPVU߉,�,V}鴹/�;�6o��m��n�7[����ɾ�����k�Ȣ�
˱M9���LvM���򪢱D��� ���G����ن��^���'��>Uu��}�~�j�@�?�nuF�6�3Q�=���G�,����������>u���~���u��^���a���凫G�@����������0��:e-�x*��oz�a��@5�Oq�23v#e���ڽ���Gj�����ɸ�ќ�.g?#�AU�h�u+���W����$[�<Ay96_�d���æ�����d�~ka_�����U7���ѵ4}�բ��JZ! �����P�,c=*Y���ޱ@ON��P]|`c���?J9�@^���f�ck	���jfz�m��\G�K�&�S���> Q���ÃG���@Էu��zag�� C�� ��'7w&9hn?/���d�紪�K����u�iĦ�$��%�sY�ܡͷ���'������E�VEQrh�E̔5���� X����6�-�ne+�T�`�q��_�O�k�u]��F�H�X�M���/�疎�8H5��ZoX4i4O�lҍ
���=��I�<ޜ��!���(f�e�j���x*�f�r�y�����\u�mQ$��6;9[�Z��ݕ�$��R��C�E�&��VMyn���8���R+ G�˔��1��y��P���$��l�u����i���elج5�*��^a4\�n��i���������f�*���8_�;�+��è�3�G�qI�A���Ў��'��m�}k-��d���#���X��Qp���<lS�a�L�}Ty'v+|%�N/�Ӧ�tf�n��xtJ+'T<o���tCXM��!t�":aB�.f��Z�g�	��u�\�}����n%8Js�=ʇ{^�7:�8��$ S�ꙏ\Dz�-[f�Ik����� �+��B��x���f2�����3λF,.�R!h��(��ݙ�5��	�yq�:{T��MJG�M&s)�18�*�z�p!�neP_�Z�/�&9T��ȼN�����Bē���	�U7���3};l-]~�6�t�|�LR�\k�]
@Q���}3��Sn�H����Z�&n��mJY�"*��=��kx�<d;I��}/Ҙ�?s�R�)���莝{ka{�;V�d�CH�_�B�/
��FH�����p=��N�17�!ͳ��\�!�%U�T`'�f\���[��Y����3&憀�E��l'9��{S~3l��q�&*8�4��6��s��'���	��V�Wޕpy�t=!/T\��
�.��G�6h����Fu��I�F[�1;��F�����_�q��b�����\�Y�/[�sf��Ѝ�U��i�Sx���H)�kG���s�,=wf8���Z���z1~:7�C���A
t0#�GMHw��Xol����ˑ]q���[��wm��ef���_��j>��� k��eF��|Y����i^��@E.}�H�ֹ+8��*��Lѐ�O�!�S�L/gl����éՖ�Y�2fa��ڍ,(�(��E��V�f��ѹ��V3�/	I�A�������L�l/�sb��ԉ'J+t��9�r>�C[6�$�W��.dk
�����tϼyf �%���<V�Bfӄ��*n��8:zf�\ར�����ulc��q�����n}ږ���5���fl���O���qQ���BD�Ó������r>z�L���h������-�@oL`���1j�؀��ͤ��}���幝z�Mj�,p�����w3.���.����rf1���+�n�\��{Ǫ*���3�\k9l���1���{�"�i0�F���de�5�(�W�ɤ�v��K�JXg�h����|u�Å�\�`�xf� ��7����A6{��M,1�s�%�j�~�Y�B���a���TWO��Z]����Q�0�|v���O@{Gum�56�����i��mY͢�������ߣ��A.D���S��e�TI�U/mf���/���A�J"�U��IO�~�M�{x��Je��tt��U7+��h��X��H�D��n��$:E�:y]��++xIm�W��� 	uN�E�ȶ:~t.����V���\�@_��,�'�������@�f�3΍մ�: x)��t���7ڿ���d�7�)���_�Fk��̆ƋT{��'�����s~/�i����]�W�W����x��_Z4#y~ԿK���Rbw2�
r�pAb
}aB�`���4q�5�ί9-E�.}^���	��U�'��n"֯�����Y��R�����ZQ26�Lhw���nO�ؿ�#��."��,�6��,��%G�<�=��wm@J]��	?.�3;�Z%u�" g~��s�n���L��US�dV��]�!�Lho�'���k��&6[�7��!ˢ�B/\ñ�C}�e���M%a
�a�}��y ������X�A*2B�y4 E����ύ�9���v��C�a���9�5y�E�c�J-ɜB0�D��ܼ �J�n��@{�F��\߯5t����&r_TZ�#����B�lE����>��|5���mpUf��YJ�٥P�U	� �S�3	�,�>��Ds�JM1�ZAkV�O�����F���B��>�P|�t�����3�<
�հ�)WB+��N#-��H��]V�7z�#���3���yAb����)��\���3���8:�r��d-�qo��0VR�����*����k�C0@=K&�zߕ嶡L����~�!��ƪ>� IJbxolk16y� ;u�O1~� ���U*
�u"��	��}�����yЩ��>^�l��R(��Υ6|6���^ݡ[({�5����k�:l�T�X
�==hM��hF��g�E���hR:�UG��C`��@w��f�hO6O�U�^"��\X��  �����w��2)#��d�7���_-�O�jN�ɪ+^#���&�HIo��+�#wE�%f8S釣܋1��P�C�xU��P�ķ=Pi�1�|"z���׃����Mv!~����N�c�1m~Q�R�r±Ic��x���������OXS�1�2��A�&H��C�%v@d`7~�[�������#�e; �
�o�Wx���#�t\�_��a�v�d8�5,�Ț?h���qm �
I)ی#����<tt��{�׭8c���	Nvg�<�m�	���ٹ��o��ڕC5ʏ9�m} *�=�h�3ՙaB�<ڃ��uRh	��kli/d��Y9[��"�Qq:��C��k��`�!������
��+T��&8��$�&���d�s��U&MÁh��?���ρ���3�D:����(��IhaJ J?0$#w�;�5�2l�
��B�S��AmR�uk�����d5N���.ni��_��I���6��b�6�1y���M��Ayr���ڻ�)"Y��K���W�X@���x��+�D���fi]�l��+����w7�NIn�.m�O�E�A�o����n��Uڕ���_�Dj6��<�G�<^jn٪tkX��p����e4\��As��fm����g�Í�Q�픟Qw�&�z������ �)D�І�v�'W�9�c.eW�% ��Œ���ѻ@� ��#��1��:�GB���II�,Є���
�֑]����X����3�>w���� Zq�����%�,7T��c�I��Y�w�4ra�qoڭ���ΉW��&�2F��?��.٫7ŋ�΁�j�C�;Ʉ�u�֒IJ�9���|i��r"{���vl��$ ÀV�C�����8�h/ni�tS=����/������dЃ`�J���5N��#%C͌Z׀�7w�G�h1��m�F�q`���o�R���
��R�����i��	�H3�S/#�Bq��0�+%��Ͼ.�}k����=���p,�D�B�Au���%���r���Ϻ�W�(����g�B���x_h���Āѡ���0���}��H�&Lࠠ��=��p@��g_���2�5��N� ��7���*GU����S�gԎ!�.�g�(8��TG,��c�U.5Z�
��i�b刾%���[ �*�������k�{VB�;A��[���2i�z" /�u��Cz#�l$��׼A�pY��Q禋��������q��(�\��|����݁�S÷��De�!�ۜ��_����2���0�\0��8�E;u��*}o1�̻C�T�e�7��(Ҟ4�i0�;2
�����s;��7B�c�u�`g��Y��(3��'ޙ������ϧ����g]��,u�3o;~� h��#|�%��t�A��
�q�m�Iyb���0Av��e3?�m={D}�捛r�0��T�������� �K*�Z/q0�fF�"�M�a]���0UJ��slQ@�]�/q![t��Κ��7i�e��-�?�rߐ��fU�W\��� AẈ���x�C�D�d�#u#H�M�%��k���q�஫��𼲮�/Ǒc�\�0G��ϙ���W�!���@���pd����x��{����TX�Zº�:�]$�d�J���\��\ U -ʢ�)M �F{=9X ���2�8���� ��H!��o�����[�V���rhCH=CcWtÒ���X+��M���.*��f!�U����ķ}W��x'd�㽲���k�Q�>�t�0XF%�!]w��
Ķ���c�[ϪF��5�67q�ׯ��`8P�:���R"��D�q��=5:���U��h�f;�s���au\��Ur?3�:pة3��-�4x����:VJ�O���'h��!KK� ����� ��| ���0�����u'�eD!��T�8����'��J���'�&�����[�f�9N�.	��j�m%C;�����9�A�Og>f� �Q���t�K_ХI���t��fK��л��5�xk�a���$�4
�Ui�:?f���$�=�&��.�cE�dJV���$꬧�NP:��%	�(2�-���`�oкl�֑0Y����`��bj9�9��co^t?4	WF{�Du��-�T�n��ZgD���
k38L���Z ��D6T%���LJ���/7t�}���5�Ȫ<=*�r9���~U%��ہ{�ݵ��'���6�K�+>�-���屎q7T�?��5`����>r��-{��[:�~��/�}M �{�ݬF�#�t."��4�@h���ێe��@��Q��(�Q\��ĸ"���t��Zj�Pމ+�.<�߽1�
�����Ǉ[=^��R��*�á�yy1D�^�נ1��ӦNSm ��w(X4SM����U	�ܚ��^H����Aŵ��(,��an4l��F$Yt��m �Qc:�h*�\���D�X}E�r�9k��'���G0~Q����i��I|���a��V�7��Hw3�^\1+b8�7��\r���@D�M:swR*���չ��_�ڱ�PY�1�=�G� x��4�*�Dg�,K�ƞ��f��n���F���de졿�[�U	���œq{�'�M�5H��?+2�^-�nv'��Vलq(������>�H�d��U�2���*Bΐ��M<1
I���!��U�۝9���]4�md�5	��ۧIi�)R8Och��&:8�(#��V[�NQ&5�LxX���> ^von��;�q�3��[�ptX�[������WNz�"�$�;{cy�c�פ3�=u$nv�r�T~;��әҪc��D�M�U:Ts�)��i��3Yχ�z\#_-�6P�>ҙ��F��alt��s+�-'�)<Ӱ��ͽs�'^�k,�P����Ɵ7ǐ�5�ɕ��`��w���
뙜�"'Ȩs���{8�+2�h��Di��C<�g��i|�>�Rw5�!�m�� lEy�%�Q��!���o0� �m�J�Z�����W��.T,���A��@��f��!	��&!Kj���m�G�AkC ���
��l���(����7A��N��Ie�F���Vc3FQ����_:�.��o,ӯ��X�-$�D�)9ǃ�ZK��ʧ�r�[~5���L�V��ꌶ�����eó������ E�)�%�l��`h����\�3�,1\ھ�;]�!�¹G�������P�٪lH�-�d�I��������S�P��^�W�]���̠���;/7��)��XsX��0�a{v� sNk�� ��Xݜ�z��}��{dxk�Y���&���)����s�C':m䄛��������3���dI���/��M��#���+��3{/��q�q˿�a��F�R��(�>��ph���/Ai9�ȳ�Yj����,��oam�_ǚ�7�+��?�K�D�R��Eoyr�l�9���o��`��`
����h,>��%�B�$ʿk��\ܤ��
��/m�g�;i�o�	1���01)���T�V2hr���5�s��)V8�]"*���%2T�7��{�:̦��Rc�X��tDH)_A�n�yX�6Cu�Z���֐lU�)�}�W-��yW?C��y	�،m��z)�~!'Ҭo��b�7�UM <�t�
9�7S�w.�|��>��,V00v
A�Ꝺ���02#gn�A��,`{����T�^��S����W29m.}^D5Y�%L)Q]+�>��.��ް7�T9��لm	�Z/&B�0�]s%�}�-Ѹ�D�
f��	Uȭ�Wݗz�XJ������,m&���j�8���E�n%]k��:o�\�U��a�\��~��ߛ��5�e��O��ӡ_E��ɋ0n��;�@t�j!쉕�RX���E�_����ӮX�nU���$��u�7�K��u��-긑�D��r�"��%���|&��C�tC��+r�#��,�h{��M���3���*&z'��s���PӨ�|k��r�,��	���s� ����e��kN�C)�[���ƋU�Ș�a�6��W�s�)�>�vK����f��jC;6�0�5����qns�),�����E�ZNw���V䐹 ���`>_|z��������}p�p"�n��k���c�׸0�#�&Wd7�w؋������Q����(n7�F�5����hN{�3v����Q���v6��6�i��Jw1ݞ��s�/)�a�N�E7oS��,Y�#]*�a�����i�U��M;����1�Ǌ��]�V�'Ɩ��$���d��h��,[	�`f<�Q�が�zk�˹d�rVr����;��M��i��1�Ey���,n#é�-r�)Z�)���@t
���F�M��?�<`D
���7�D9$�6[�k	𧆢3�]��x�)8I���fA�G���\{(q���Чk<-��!!��>g��N�

)�\��Z�6�����.��| eM�^��vQ|��:
a=<{˸X<��5g)�z���o��e�N�����f
!�*շ��m
p�"d>Ui�[�~�n#�X���[!"�����	������fJ�K��jě�E�6��ɿ����������Ԋ��k��;V"��0��T~�ض��Ib�K�X�"���]��˺��FF_X�-#-,�����{�rS�|<�m5IK� �9.t�!O�*�T�!� �;2�F��j�N�H�j�/y�{���������5NZ�8zÇ�;���J�(��8��
6�z�'Ӆ�#,�����?F#c'�����E�J���DU�L{Ct/�Z\���	:�Ȩ��S����1h�]3�Tq��Y��Ն��)U���N����@g;oa)/�}���*[�U�� ������"�3�i��vv9�t�� �R*,�_���ц��#8,��m�e���� �Qt��^�SБ�x�O�⧆��II��ʝ8�`1'&U�����k��Aֶu�!�m0����
��|���Fo��\�m�^��kxC����Џ;���=��
#�)D6��CBE�U�갮�.�P9����lAX4z�_jt�N�U� �l����0uY��c#1:�B�>�Sw���?N|�PX���*�u�3v�,aS�v+"�j�w�ϲKP�hk���ôK&���WM2�j��9���1�|�)uk=4�5�_��D1F�D���J�5}L��s��"{X��xu���e�`�=񇱳��+d�2�w8-Z��j�����pO��&�5�>WIC��D����޸gu�'m�sjck�; CJ�U���(�g$�����e����Q|�ĕ󶑢�E	�Z�E��%��l�,���F��/xjz`��?oY�G8ҥv==��������bnLd��g���x/�N���]{)/���vZH?>Ee�I�/O]]�,>~C�_�; ���6p@R��p�k���z	��ltp����:7߳��α����b���j��sY۽;�h��_DC�!UAAi��},I�Q4=���&G�2�i��}Q\"��R��2�˷|LF6�Laf>�3A�Y���Hei\O3���W5�3�ƨ��`hU�W��������ܞ��;/M���g[����,��Y�	f.Y������7ׅ[��HI�S��s�#�A֝�"�7����(֍�4����q$8��i==K��B.�2-ao�A� ��*�YGr���޾����'�*f��;��)j��C��mS�X	P�>ެ�Y�Zw��G�F�R��<v�)]c��ʹ�����Db�:*��FK~���85�Y���'[���kg�;�
��6�q��]7�
C*�B����@�t��C��o�@�
��p|���j� Ȓ2D�p2%i�\MZ����~X�ƭ�oE�����g�pJ�J��8ˇ�B��q�8�Y����;$c�k�8�"G�������nτw�ٜ�e�g�2���g�ڕZ��*U���=1{�>�˶��zك�t2x��������ݽVi
��_�4_�~X���/��p��ð��s%���jS�o��qZ	��}�d����軥m����N0ǖYߗ��A�h�w�!2�R��ʠT���A0��zE����N7j7�����`��(�$�Tf|�4_̚o��.�������i�P�pR<��p��2���7�(<!����mb�?ײ�s�n�Q*0���s����.H"Z��b�#ӡ����F�FO�v��L*-�xQ������q��5�:���HUnǶ���=���J�}xt�/1:�:?P� ��9}�{�awB�1tt<c�l����7�Qe�+��Gan���x͆&>�]6t!|[��0�y��ԣC��$�$<L��a�aL�Ϳ����^�p�~��Dl͊�:��枈*d���\*bM�BN�*کݔJ�\�@Ƭ�c
���;�������+Xr�����Uq��paB�����@4&"�c�1���D�VS�6Å]�$��T��c�c
�s@�4j�̈s�Gs�\��qZ��TrÖ�n|x�OW#��aUg�rsFi�q��h�����F����%
�)'&/���;�Vý�:h
��W�Cgf���3��N`nfkD���8�Н�k]]�a_c5��؄��5��)�b2�8�G�,}��T$a�'��^�i����f7x�8T��&�;*�_�S�Z��\�tSp�g���q����e�P�ݫm��R��ߚ~)jgS�Z<�^�/��J4jR���0��1��y��ΐj�@=Z�V���'��s��8k �`��i;��8s�� mx��F�RWFf�S�I�� ��2=HqNBqS�
X��Tw؅� E+�u�dI��Y`"k϶���u�/0���\PV)vJ2�QY���x'M��ط/��2}��Ӛ��g(E��~���hh�uJ���a��=\\�8�A�[I�n�w���,-#�>2� R��bqdj�$��OˬH
�n�� �j�>��hNL/�4��&S���*���<�s���s.t��[aN�Q-`���3��n~�M��e�:)��f�DcmF����3�3O�
���^��\�)��+[�'����.fnw�;�oET�cW������d7���k԰�a��c~��Bo�HuB����Lf~�ܱ?��6��E�,7�C��< ��9������j;R�HAD��t�jW�a�1�(��ي9p�cl2I��)Z���r�FSI��ԙo�nw�&��Fh�׶��%�-T�4#�ܶL8(�yՑ�O�fq ��c�{�?�](B�V�&�O��L���� �g�Kz��}�eeA��8��݌��C���UU�w�d��l�X<
6N?� ���	�ڈ���U��N�n//��88%~c�=o�=e|���,����x����"[vP�@QǦ��E��`�!�ʣڐ
>������ ՠ�i�0UU�D�I�X|�C��5�;�׉�o�T"e�9��6���uXV����*xcs�z�:�O��b1��C΁�Oɋ�C��J�����m��p@����?;����ɇ�J�'�M�n�g��Mg���Bj9�P�grlK��"ϼ��j�Sk8˫��7��/@�R%d�����g�3ָ,,��)4��L��f�����@MpI�Kk��/
?�LV��/��m�!��_�+��:m}�H<c�h�->�/�L��>q�6s�fŮ��Q l �NL�pr3�Vn������mv�ԇ�&$x���%jD��n�-�)�ޖ�z�Bfl4�v6j��ԡY�AI�����L\Ƨdӡ@74�S�0��$=���f��b��x��-2�Y������ofJ����Ab!��<���f䷋T��'���t�G%;AC.uB���<)n�eeWnV�A,�ocX%�^�&��p�<�d�qXk��`�S̯k6�Vٝ�����Z��E视�̽�ց��*3�V��c�?6���1���H���ZTe��O����Q0%g���ٰ0���Qi�nc�F�ǣ��S���-Rc�v�͐�z
̂��`L#!~TJ�� ק֎Ӌ!���[�1����Bs�| ��j��B�x/�7Z;�9ܳ[(X�á3�;��3w��}Xѱ�[㜜�����6�{'��WO�ÈT��\D���<\c�>2ڕ��e �V#�~�h^pN�т��Iwj��]@����f��OT'u��56���P!��N���	¯�E#qEYI`X�5
��tbA�s�_��Z�e�|�`ǅY�����68����e�DOO7MMx�!��2�i������}�@�� 3��`Y��8Q��Ż���@���Eރ���	�O�����̀�.l�2a�þ�~�V��������y?o���,���X_�|ﱩi��E\^'8W��D�I���cXI�R;�4�)�^�Y��0����H�?)��r9r��~X&����K1jt��$��$�?���3д�,�R)pFB�).2͠7�%]!�C���c�B�3z�N���	��iŨm6?�q�|�:<�9O�=����[�r�6ӆ������T�^t�?�Iw+D3o 5�,�r�d�d���| ��g��/Í�� ���҇�����F_�[���l|)x�.�������0�s~�UI2��L�x+����p Js�5����Z�|��n�3�:N�d��2TͶ��K'[��v����ee�9�&�HY6���Qȱ�<P��/$����n�V1�~���K��:�R����V勯�"�=�ߨb������;�Nm5��״3L��6
�}��`og�4�n2Wm��:�ٗ�?��6Ji�y�7�Q������2��L��@�aO�����Mg?�[���L�!�@��+}O< �=�;��,�TG�j�1�|�jP��ı�=�5�#�����M|�Q���/N����A�ga�N�^	��	���Y=��ٵq�m��M=��Ȳ��o��[$�-�!��$ÁͦU���ݏm��![k-�
Cz��5|&�����4�$�q�ŝ�i���a�Qk�����
^}>�!��m������v_���qf��M���`H���I>Jsf��K�{>�a���upE�#`���JlT>�X��e��xM��`�M0���ޫk/��{9c�w��K̩B-s��Lp��J��b�A����>���h+�3��U�d�w�%��:��- �6#��l��{�j�B-�  ������F`NP�Br�f����g��O�Qxa�q^[�!�.�1�c�q��8y�u�&���~�?��Ÿ����ȑVp��/S�|��)�)�9D����Y5�|ߝ�1��ÿʶ6m�Ӹ!���G��!du��k�c��w����uD|�P	��Y%[����+�&+���TCj�Ua�ޝ��;�0:ͣ8�	�w��.:#��8�Cch�l��G�I�d��Ck����2�5��O�����BQy�6+Q�A0�ҷzlԴ׀uM��0_F�FJ���$^��ӣ�&�P�Ì�bԖ=�T�2�Y­6��*�%�.�gb�Ϟ����7�";n@���8	S.F<�""�y��X�w����|��<~t�<��?D;�V��ݝh,���p� D��-]?v22��X�a��w|��:f�vn0^������	���_��=oOyg��ԧCaP;�}g������9�
F�"�;^[���'y$���m�,��V�W��p���\�C�c�����\<[�_�=~. �k�Θ@�I�TϚ�1����T��N�v�!���;��қ�\�x���֯ ��Kƻ	u9:��� �B�5z��Dq�_���&�2�y(_���N�!�������N8j�}U�9˹��6�5:��F�S!B���~��s�03�M����cnTG;�݌W$�9���nU[[Ҷ �����B6Ҿ�p�n�>�VX�=-�f�t��
�F�kaHڙC����$��������=h�������g��)ZY��y��]|����Y=ݦM�検����յ]���"�_=��.Ӹ�E�<��)C;�6� � &��seIv61�loy�,	B��Gs;M��f���,V��?�&�V�0|�p��f�^[�+���(�]��RäC[����/n�����_�N
�� 3�U/�|y��hUf��e��ֆ
���qa.�@�P^$|(�碶�W�X�0�_�W���9�ʏ��X����0�}8�Vz�;S��d�[֓�9����8�
���Ȇ�:ڧ���a
Oj�NU����/�߉.�Q��2��h��T{^-�	n���|칞�?���^Ӿ�t���RYt�~��s�t�p�:�z<��}��1_2����IM�#�6����iRfu�}�'���ZQp&�7j�^+�S�?t����Ł5f���f[����w��Gg�r'Q܁4��苈)HǶ��"x��͆�0�Ǔ����L�o��}36]gK�4^�N�����蝿?��u�+jy��!��.��!�B�A��,ʿ�fɹ�8��r�mrNd������Sݽ;�\�,`�%N|/9�=տ���=�h(=���^kg�M�&�C���f�Q��攔�/{i��C�]~�m�����eT�|�Ib�S	� �mk��B^ɲ��u�S%�$nA�:�5��m�Yy[$>�v%O"��с_�����ڣ�=�{R��������q|+C�F�p�F4����h��AxNS����1cE�5�.r1 ��7��0�2J�	ͯ����'R�h-(�_C;b_S�(���~H����w3�,�5Y�f��qS�V���xi��IB&��_6D��׈��qv��E�!���Q�Bm"E�K����!����G�Лr�'��눌4`����Kb� ͘�Sȴ�S������e��Y,h��%�=mçsZ��(�w�p%o�8cc� s~����}t� �Fa�Nߑ�h#Ӥ�!n���2J %�Q��D�aV(:S+���L����r_g|o^�a�|��ҁn�7��*��E
��cJ�i;���3܅�f�{If\���-D�h]��N�Q5ǟZ�D�ӻU7����`Z���:��t�!��B��a7�*~A�0���@��2��C���*�5���i��5~u�9yE0�mZ5/�P�����=C�L��M3�<�C��iԾ��?��;.����ǒ�������'lC�´u ��-n��@��!�|��#v��
�;�����Ʉ:ƺƜ�(�lA�% ���C
�2��7wl:���c&�	IߨB��C���l�����$��fUZȉ�	�R./2,V��	�������\�2\_<s�����ޥ/\(x�򜚞h�׊<���]B�D��꓉at;A����*F?���Pl!��W�dDc�o����q���s�h��H�V�}����#�@M�ݠ��3�qkGF���y��o�-H��h�*}�F$-t�W���&���S(t�(���绉&iis�Ҭ��I׺y�&�C{0�8p���2��R�	>ծ1;$C{��Σ�^�p���:8OJ!��Ϟ��?^Y_�;���C��W�Ǩ�o��Z�R~w����nI��&�_\V�+y�#�D�����f���v����:`����%z(/}�<�gu��i#7���Ĭ� s�
\#.���;Q�O9p��[�= p���y3��K�Θ��(��Q:�c��5��h*M����]�y-����SG�b>�6;��T��Š�mc�']�*~&���S�����	�|9�75���}��d�BE�z�C������d�y���K���b�-`���GO+�N�I��/���?�kc(i����Mu���}�#���z(h�e���mh�gr޽��2�[��0�`BM��à{�7���d�~v�6�#h�ҟ#T���8�6��1�m�&*1a�r���W���<��`��:�e�9�H��)�>�r�$���V�SMz�X�;��Vj;80���u"��hP��2ԛ��vF�-�;x̌�=(ǥ��/����]��'���0�����샜JQCu�6�e�>���'��}(t�\�p�/���O�}H!T�<�U��'��W���;M?��&�b�!p�i��gy�<�HP:�CZ:��}�o|��>�"�AˎF��Bx��������i�M��#������z�io�U�ؕy# ���-C\��fg�B�F/��H��B����!S�a��ۚ��_�w��~��'�7<��bv���G��(Աf;�;�w��|͑l�A�����?�[���8)�b�����U�-�#��:RGj���>�>='��{䁖�ybW?�:�b
U~�{p���R!d���Rm����Ι�r9�(W�)��Sޥ཮����Y*�����>-���T86��F2�kZ+�lR
��a��X*dN�U<�p}�y�p�z�k~�Lx�oI���a�����Pl�3#ዦ�H�r��-��4�!��T}f��m]�;��!�ȁ�l��K�'̓�iw���z��h&�o������nֈў`�9+��z�K�5��ͅm��u����d¤���?�ZK �<�Vֶ��&��`� �K�Ô<a�=p�޶�ۏ�9��{�Tu��i�]��w���a�XYZ�z�tl���MQ�ύ&#�,��A��x)���;����G��#G����ɹ�n��&���hQ�)1�����<[�7's��=��I�@���}J�@��~Q�`�x��X��s�6�-��C�A/:�60��H�-x^gu~�z��5��8Q���?�M
��p�*���95w����,��; �_��7���Ҳ8�/"��S��*��p��]�6�W�*�����(�8�D��Yf9��`�J���OV�ְɳ]a8)�s5�DS�c�ɔH��f֦J^�h���qQ�X�&��Z�Cy��I�Y��.�ʺ�كe���BL���>Jةh�j<+
H4@<T)Nfz�GOWb�qL�1֡xe���/�d=���b�+�_�E�I�����Is�\(*�A�0v�^�jLLA;�<qh��ϕ��!�)���<P$X�!�s��`em]}�рڜ��߮=��f���}��H 戂���r�mn��݋]��݇8�U�����A/XčA�`D�f3 /X�0R��Wn�V�7�4���e����ۮE�:�oC���>~ʰ5��$ÓO�4�dm�/IuJc�����%ߵ������|1�����)E*(��|�$J�p4e��#� �TeD��mI)E�܆�}��0�QM��=/\�Qk3���*4�?vC-wW���<��D�'O:&[��a]9�i��tۥ8�_q߁���]��4��I��Lq�|E�.�;B������>B�� ���/�c��Z"c���fZ�����K˶�|p7��؄1�������w*$�S}�!˙v�e4k���P^I[�Ŷ��-�>!�ٓ�F�Ǥ�c�1��i1�[�a�Z)���t��J���c�v�w��u9%[F~gB���=���9��9�sv��9Ʋҳi����LH�H�.��';��P�Y'h;�l7V�������^N�	yX�+ё[��r[NsGY�6���9�i�%{�q�{L���ѝ�X��Kx1�����Lm�Q���S�(���lPVa,m�lrFB0�\om��,�$�3�M�eqh�K�ٓ_<mRp�Y�QCFl��߰}ё3]�.�x���E؊J�Oqʳ*��.��!�KC8�ʨ���/��q�vE�`?@#��I���/�g�qP���FԽ��C�0ޝGrϿ���q>���>¦�O�
�a3R���j��+�T1�K��	n��pΩ3��NC��I؄&�7o�$L����������n���Au�}y�����p�����s�Y�`�(_�z���6/-f���Tw����ik��oY������Daa��x~�{�LfG�lʥ�_Q`˩0N�����;��r��H���)�*Z)�I��`���������Cdlc��2���ߺ����(�������դ�R��f�WU�����L�{��?'Lx�C4���ł�Fl��A/�6�?/W��fN���f�8�m%&y~`�C{���T��yN��E_6ÉC�.ϒ�`�U�)���/����~�ɼ2�	��(`���EC�48l��0R����4㶏���Cx�O.RM��S¶�\-��
5l=!�G�B7�xDs����`�����͵��7}pZ]�.�#�DO���	��,R�%�*���A��tj4U8��"��FG[~m�v��!�gZ��Ȗ��21�x�]�@�(עL�v%����&�3{+gj��x��q;Fjj���M|d.���cn��Z��_�0A�8A���jw�ծ�󗱹Qe �2�����vc[�D�>a��E����Ҙ����q]Z �!Hm�W���'�#�`����O��Ef��Abox!�m���e���=�H����	�7�7r��K%�p�z������a�mAG �4~�ޣh��)��J0�H��(03�)i��PŲO5c$Q��O���܌v�5��ƾ�K�u���*�d�C~d��/�Yȝ5�^��B�.������jq���A���B:�_Z҈'
��	�N@)K��?+�9�$$�4�B� ���yr�vD�Gh��@
d����v��r!�Ghy��\[�X�Ϯ������*�\�O)�A��[�o;�V�c�x��}��I��������v�w�\���z�_UV����P�A�|!=�8�Ur�l�m���B2[�%b1
�<7t���o�m�G��?�kA�Kn�6��Y@x?��~ؠ^�KqL�0h�K2������[����xF2�o��#���"/@ԛ��wg�o�CM����½��O�$�UL[N�y0V"Q�p�z��rS߄��`7�2�ډ��ޣ�
����+R�,亇ؗeMz��s�K�j3{\`Z�ps~q[����[������X)u$-G��H��c��K��E>�� �j��GǯS��B@��9��<4߸��(Л�ZL����`��Nq��\�\׿�H3�A�v��"*1��\fJa��U�;��#B�@��Q�5;�bJ�p+ºj9��T�T��*c�HA��l���vHp�SK����uf�u���;�����]�1��n��M��H�\d������h?c��F	#�wH=n=�+�N,���&�����;P@��ԹDW8�+VΖ�IQ
�m��8����D�f���j�����O���+��x��f�-x�ktȻ(Ү�,�=6T�Ǎ�1����f�.��p#;��5R��"��=.p�N�Ն1�8�N9�F��
���C�X��u��y�xV�2�-���nQ �����!�´3�4��/�2���#w0��v<�������Qr��b#�ޤ`��EK2ƚ�F
�t��HD� �3�Q��Jr�� �L1Ю�W-�e'rU�l�f�����<�D�}��o��p �f|A��eG�ȃ�n��)���6�^�,S�\�6�7�~QX;z��b6Ơ�kM��c����ɠ�`���&.�F�����>��=v�U�!O�8{��&E��&i�>�*�u��6ޘU)�qWG��y�$Ԗ�|�(�S����.=l��rd&�ka�[*X`PJ�,c�e�}`������h�R�P逝5�uU�������#ώ;'A]x���Ǭ>١9�i�����%��4D�S�	�VΝ_�S���@֊���k�[�|�C� 7�!��n,2L#�ՁhQ��,L�>������c܀8�	�6�a0,QĐ�u���A��Ȼ4�	���oҪ��!�%4��0!�B�n
�&@��9ob��	z'�-����b���	ĕ3�LW� đ�!��ӣ�i17�
�4*f8N,�]W�3���H��$�!;qJ�F�����I1�P�m�Q9d�p`+�o[�ZU)Q��9�kʫy*��Ww��@���eo<�9*���R����µ���_wV�vAJ�"�.6�������og�m�,� �*%���Bό�KC���_�����SA��~\���;)9j<K�n2#q���)��f-@�Aۭ�v㒑�P Xq�����<��ө"|��ѻ0pn{�3���/a�>r��Cbjo�����h'��:�_�d(��uF�?�Ќ���<f
+�#g��$"�cD
5R:aƋ=��t��I3�F"C(gA)1Hr�X4vZ���Zy[�>���Ð�"N!td��c�`
ro�aR��y�U���o%�1H�ۄf'~��<�E��7[\������������3g�`�-�j1�-��~��.\����k�Zh�G݀cӣ�8(�>��h���QB�I�< �.�|]$AG=�1��8r��C����<�,�BL�hO���@�a����m�	���٦#�Aw͢�<�f���Oc,��ͨ��(����4�`����w|�c�C��A(͏x	D	'T�d�Cܾ
�NK���U g��雈k@�|��H�w@�Nk,�IJ�GԌ��Y�RY�a�-԰�	���HQ���_���`z�D�y�����yr� �2����1J�c�2��J��M|*Ovt.)��P?w�.(J�wc����� +��Q'�����i}O���x]�h򙯦1O�2嫫��*��z{�o�:
|fkZ��B�=�2,,�X��Ms�,��̎($ԕ�P�ȼX��;C���rh��y�E���sߏB��D _4	 ����Ћ-��M�x�Zʤ�C���*�?�M�w�Oe����y�~Aʚ��W�D��2C9��Q��87��C���y{��mO�_��l�wJf�2��S�y*��f\�H݋�5F�u���lǭ_:�u+�M��U��UX����.Y�F�<<�MKC�{��/s�~<� �J��3�����������rm��A%7g�n.#�1N�@e�{ݩ� f��|L+碡K�V=k�2�b�s����A�sEb���%�2Ɲ?�v�[,?�Q���	�����"H�1���R/�}��IF�&����hQ�Y���5S"�{�˶�i�]I�z��s&������k��\���ƔS����Qh��k�+����w���wb��&Du��O"�	炩F���Ɨֱ@���fgDo@��[�d���$ى�(�p����ʾ�a�Έ����N���"u:2� �D�ۤ���7.!D�-������JGo$����m��Z����$��δ�:T�gi>�#p7������)� �����c�w9���?z�4�8���r�҆����fp`q���&�af_#��G7ʾ�j���)c���a�,��gJY���6�ȵ��Tټ
��T�$�E&i��y���f��*U�0�{N�����z�x��s��Հ�v�P������m��4
ƔMH\��[���Vh�!}��oB?�N1�&ͱl<%~�f�Z�YV�Uڰ�c#�v�bFZ���[b!�n�t\#�Y��~2�e����,H�~Y���6G'�Y�o�U��+����!�Za�h�3���MV0尞u˄��e5�Gv.��Q>X��]�*D��\)��կ��p�
��1i�̉�Um�'��x7�s��9�Y	���<��i���j89���3�j��r����6�N���F����w�m�wd��|�Ҿ�D5�ekx��y�,o��p~j��C��kj9 ��HGX�����|{6YO�)!�w����W�l��������%k��F?������B'�F,�S��ҞU����@��]�W��މǮ��H��v*%@����3io�QCݷ�D0�7Y��']��y}��ZB؏��?~v�(+����+(< ���}r�8��_���7L5��9~���gD2�v��I�(��l+�r7�e�(���P���[�mZٔK>�*rB|����k��1M��������Pze����5%w�Ogw���ņ�6E�z|aP$�銭�� �F���qЋF�}̑��R�u���&�8q�$��o����l����|X�%�C��{I��fgzCE���v�h�����{`�+�L��L+��@�ʟw�K���Cl�*_J2s�,�w�e��w�����c���yTo��aBYvP(�[�;��mM\��7��';2K���'���%��h�PvS���Ս�b�7%x�?i���Զ,������:C'OT�Х�'��MAEm<:߹?M�����oF#�zǔx͏�Q+k�)K����È<��6[��H�R��\��-�h��~�C�QX�r殼\ή�����Ay�i�*'X���\�at;!W��Q&H��y����I��mۆ�8x%$`��2����Iܪr<��*������Ajfɘ�'D�޻+핒xxO{g���H7K0[�_�zT���k�����*E��G���T�����+��<�)B
�S��t��h��_� ?]:�2`�wS��435Ρcp)O<l�9�`to�K��ݢ]�aO��h��d�� �W�����U&i#�z�����x-h/ �_��IRr�>͕T�!:A��V�'�_��`�/¼�v
�����UR˂ru�-\%'���5)��؟'�EƄ�4��v
G�D�%?4��!��0v��ݲk+��a�Zo�~��� �݅�I�?A4������>�fݺl����`g�2�u�@��;�*ɂ8�N{���$��~��<}Iޝ�]�fZ�7k1v�L؍w�U3JWHڎ��>�N}�9�/$�F�E�뾴~��1�h�3��F�����mQ;��h�|���J�Г&�s�&��q� �HR�&��Dl����:����4�\����m8��+�P
T�x�o�d�Y�'q��4zl ��i�ZJ��</�~N�H�l���e��0�(����iA$t���$��!#�[��G����}>r�^ľdϑ�M�Na}� ��؈,mQ�JƟ��e�g��b�C�(KT��H��"�֩�CS�?�
��|���_	WR���O��նK��:����N8σ�H��=��u98�����)�ohf]�Tv�
���= ;��Ip�<����{��*'9k���i�B���5�{�7�w	�~[��'������gّ�Ԟ_t([pLXbD���4+g����~�:�L��\G����]<��� #��υ�'XC/�B��u�ϊ��
�k��܊�/�P��F���
V�-��@z#�FzY� ��@$O������q$�+MZbx@R���Q�"f�w���륩�S�"n0І��藇N�+�v�����b%��	�(�/EL�x�Ť�JP�4�"2-��#?5G��G:��64�Z�f��=)ґ���K곅$��@b45���V��-ˢ�C�V�P]���Z�0'�?�(����VJ��to1��^w�ؑ˓Yz�h�l �%E`CL���l����!����IC�[���zY(��?03P��&�����������e��0���e���w��n��RG�\��c���3��*�_z�Gu�,��=+@��~|���[������D,�C���31�е�����e'�kbr+��7���8ZJ����a�a����LB<V�}UT��詈%	�l*Z��=G
�wOe�V�[�]bj�8���Y}��W4�]| �)Px�G�7��vzI�H�|��Gf��"*�E�Zz��E�5��ژh�붝���E��d&`"�z�����|�d>�1uBHWft��������F%�*��R;�� �U݈�|��G��}i�sy�D�ɂ������-ޠ�=�}��t75�H}�[ 8�k|�`�����F�%(*��C<2HH�EN�3T��x)��;����\^�L�V*_\��E��<������V��$N}����/4N�mTj�"5MNc�U��O�F~l���Sm�Ih*	�dQ}nC�`�%� mE��U�zK�+���R�(貰����|�|���{"�M!�*����M�9�u�����#�~��ĭz�K���8d�ʾ�d6����zץl�ѻ��&�Q�6ao��c^J�|���PS�:��o�'�T�Lq�-��<a�z�x �=n�����*	��_��i�rh@
�4c����♧���t�yUۦ��D.9W]?t~��y��\�[KΑ��FI�i�j�}6��q��Ӆb< �t�Hq�'�����3��H6�ϛ�������t�ʍ��,����47L�W'�M4�e��6�m��K��������{"�7ǜ͞��٦9ml�(�E��<�������3�܆h2kO�y`)��>�OkWG�_y�8�@��F���5&����1y�('���x�M%T^��X8�CMsp�q�/w�C���9���G�����$�� /� ��Ȃ���*�2��@
��#)�&m�sl��{U�O��-����&�t��vjݧ�sDf_$��'h��z2]k��FA�o� 7��e��1a�G=��#�?�=O�s4<3YR�E�tmC�Q@��8�����0
���5
�#4����4L�|6�X�xo���=c�P~���Q�\�$$}�,��(�z�5V4.%��t�0f�|�]T�i-��Aυd6J�2CT���G! {PA����k���A��͞�P5��>�2V7�7p���-wX�=�$�����pyE]��f},����s�2�6��sZ3ۘ�<�҆�6x%`����/(Ƈ���S4��ҭ�H
�z�|��h�0�1:��3��TwJ�;�tW�l[�wٖJ��e�)D�����x���y^�2�<�Z��fW�}K#�UN���a 1-}H�N�c�u��\�D�>����=�M:��Wg�0%�A�Ɇ�h4�s���k��mS)���Z6�����q�V���4��6���ƒ_{RU=��nk���b�i�xcx��[�헠��D���������Uu��T�њwm���Ȩ�gR T�Y>}�¼��u��zBj:�'�ӫ#��R��豑����N��R͛���������fT��1�	Xr~�k��iq�l�X��(�ꃕ��T9Zy�&dpŝ�%\���_�E� �Q6�ıl�u�PZ`dr��r�O�0��&N/����%�L��@!��
[˿�?�R����A�.���&���[��[%����;J;�_��?�<�Md�n�r�#."�_=�.d��QX�x���q��P\����@-*ɲ���_��I�hzh$�����s%84L���Ϩn3T�\��X-p}jo�Cj��k�-����-D�?-��)ԧ�
Je�\�Z���Aj9:䖕0�G=�h@JI� ����.�^Y����n���G7A3�ĸ���!̺L�Ƴ���`|5����L~A�>eَ�q�����΀�e�H5�6�v��a��SGE�f���+��vۍ����G��rC��YL����y�ҐKMm:C[����Ha`i��+;<�A��P']jC_Q d�=WB<�J9v�v���hM$ �(�P�� WksWm{dԏ���%~��B��+y�L��l�d�=�,���H��'���e*�E���Z���Qw��}P���]��B��6�&ᲁn���>�y�y��B�D~'1��J�s��2�oR���G��->O��b�_��2��]�W�{�����y��\��7����)�'J�w��n։���>�q�G/�]��h<��q{3�E;x��y2%�&^�V��\3�d�W^̛؁��*��N��t\�c5�Et�Y�-�K¢���.Y��h>M�������:<!�����f�Z����G<g#@��rj(Od�'E�5����6m�����zG{=��+��X�"�� dc�Oa!M��pJ�D��RБ3�J��+Z��A���Q0]��������Zx(��a"�C0�LM�����ֻ~tM���Ɓ �JF0a�~�lR@M�1��,��;R®%��F:�@)��B��ইt�lqZQ!���R�8����K���M��
�|W@T��3�J�ZIl��5�<z�bP�/[�ˢ�;!���s�m�$V���E=P�@��ޝ�Z�H��ҙz?iΎG�XN��~ɨO�'}����A�5+d��K���gG��B(��i�Aھf��3�Q���10�p�YA
P��̐�H���i�	Y²�M#rU�u� �S|��q������e�n�uO�u�M��®&[c ^.��\O������m���f�KF��parO�p���H̊2f%�6��c�т���J~%���uH��^��G����,�0PGL[��_>��>�! ��Dn���:&	ZhRe��}�Ko�c,X������=���F�1{ »U�_��f-4?cSea�r⢹����~| ْ>d滳=��7�҇���k�s��%��b+��G#	uI2��h�UAQ#�R�[G�3h����QJ�,\)���`3���8���/ܶ�2��$�_u����a.�p�y3�&L-�̘��5�U�[����l�����g�w�I�MMqN��g$�;3�F��V��M����RT2�F�@�����j��-��&�S�L�h_}6�m��!��֍����	���xt�b�y�	l����8$W amc��D4qk�p��Z��:���������=2IpHQ��u@�_�$ۨ]E��]OL��Լ7*G�᫙�E� T�,9���.՗ �՞aZ�`h̜��:���o;�OXiQ��Y�E�SL��Ҙ%�U��,G��`)��-��JQ�W��~�����;:{�d�ʂ��C e�*��;�����^s{>��H�����!(ϭ=j�>�f4��Z��Ç�I\�/��"HW�om4&S�CK�n&�h��u�M�hYP���OB<G�����(���ܟZ�v�|�J9�׊hJ��A��6�/$!BB���r�OI���Ѹ���$.�<4�T�C��&�*�����;���"������_��H�.)���icZ�R9�)�cp@q�l�%m�|���x���W�=;��?�@,�q�=�>S#4�ZMt�&�Fs�����v�ܐYx��l������tD&@yՂ�]����D�	,����;�����b�F*��ݑ_eu���*�f���	��$�ݵ1$,�h���c�`�A�מ�y ���\p86H�~OֳKt��SC �5^ѧ݈v�|-ۼ�*0�T�;S	K�:_]h��i����������m��|�wE��nС����.��{;e*a�@)Ju�B�����q�J�FyY�ƨ��;�8L��N���J4:��^,)m�u���s�z�k���xytD����L{�-�e"[\	��w�@N�e�f�@R-��E���Z��6�,��4��`QEB��>Pc��މ�!���)g���gM�'�UF�@ҵ��{Y}c�����M��ļn�94��˦v��X���p_Zc'[O�e���a@��3R�?�e/R݇�.xX�`l��D	X���4�I�_��W�#Ѯ�rQ��� ��n���T�{���ӫ���*Ax�Tv�[�,e`<����c1�Y��T8K�>��8h�ٙȋ�\~ߞ;O�����D=ŧh>�e݅�F�5\�8J:�_�^a�Oax2iDo*草)�>����,��e5��Î(���!���|N��RݹV(��5�/�3��/1�3�h�U�������0��ԏTB[��Վ��0'�g��d?��8e6eN8�����Tm_�j
%��N���<�(���d<��q3�χ���"�ô�F�F^47��~��<����h�r��(�ܰwg��Ή�la�%�f@M3]��$y���ю�W��#u'���L�+ѣd\�.ю�r9c�]�J�`�R�;��ᙲ`Sͼx�0ntO�e<�� �%����A��\R���	��2�S�oJ �Cr�����Ub	���Y-_q��_�Lg�݀.�]����E��+��zr�d,�I������w�k�ٺ̝�	(hq�Tq7��>w���W�`WxҢ�9��l��qr�� �C����/L��>\��lYn�	GɊ�f����1B�Տj�p��� >I�ʯ�Q0Ca֩l��������b�X�}�U�S�S1�͌�r�}#�� Uj��b\��mj/��N�Z9�Y�PU�V*���L��Ţ�A�?��L($%zu:N/m/l��7�7&WL��^�,��u�%ףm��(����{v`C���X��_lWn�܊i�z^շ��wv|FeF��;qa��&�{v��D�~�i�i^F�|m�:'�	�_Thq��t��5�^��y����t��l�86U˕[�/	R.E�:u2+r�<���U-�gěkM��K�5�R�`n�8�[]]�.���2��ţ����W�� ��p�U��*�OY_?���9�jNoQ=����[�	C�}}2�N���kʳi*��J1:�l]�T�� �q��F��&�B�׃�ZJC�/N�"Y�l�����
iD���
!�z�b:��u;E����)�Rև5�/d�bH|u����$"6L��u4������s�#��< ��b���;��4D��c(�V��쳪[��R�Z�"�L���b�V�B�:�x>��;��%6Ё�5��Z�Fv�V��(�+��=Kc����B7����y���j�jɊ*,R:�zk�9�u;^�_���E�s�<����-\ߺ�d!/�Fh�`�IG(:�G��H���IG�6mЋ�P�����wۄ�j65m�#����(P@�6ϵ��\ؽ���ݕS���c.cT~7� m�b�1����{2��-d��AB
���D��hj�јT�뜻��# ���vU����Eys�������-���@�Oѓt��~`��,��R��j|Y�D̮>��Ŧ�.�+T�dܡ+@�+D�����g�|y/��g��/�[AN��8W��&��j��=lS؈Exin$��;㉙\�{Oi���!�y���T�>r���D��m4�A.:�{W������.��3�<I	�,
s;Y+sP�_���q�#�9?�'�m
�ac�'�-�(�NZ�J1��;U��������[W�fG�|���ؓNS��^�J���џ��ӽ��E%P��ϝg-�9q�5f_��-<�	�c�����Ď�e��`%8��趪�t�#���]��^�I��+�?s�3�!������%>+]+�Ho@�F74i,��o���isH�A:��8�), ��:�j�%�e��ۻ��CJ����q���4�����
�Ϥ���b�,W̹����)@-�kx�oq+qd��2�M1�,`��&��6`Axb���ut+��+c�H.�gg¾"���Z�S`C.�5yHu	���f�<.@����TG���jH1��9���{����ԉ��Ulx��Z�/�>N��I8qU�\!�D���Jk��!dq�� (E
��y��߹�Xc��G��F�S��<���〙~����j�o�N�P[>��ySgp�U�PD�#X
���s�����]䈜��Av>P�^�y����ċ�=x=CM���>ݬ�������8 J�"�>c%����ć����J���r�O��DP|g7����QU,n���)�_2�ɣ���� y��f��#+����V)5�u~�Py����͌Ų�
O��-66�
�#^�Z~��JZY��3��k���i$��A1�i������%���fnE3�kA�����Lr5;�.������{x��F3yǒ�>Ush�~��gA�^3[�㒏>!rUc��!���x�m�lB�����8��U0������h���Q���/�u�_i���K�xʀ$Y���C6�[�!�F��a����-���)>X�*ihs�����^u"����}ٿ{VP����|�\��S�c5��W�a�(���i��Ҝ��"@�T����z�c9#���p�/�����)��`3�m�+x��l+��}y���E��{����Oys�6�7�^�ē�ڃ�|Z+JM��;�ʯX-��@�P�A<����'��e�����Naܗa,���'2�Xi>�o��<[N�bδ�]w�m�A�)��lž����#1�N�_]:�Nt_�p,��&>]:Uww�͓�������>O);"��Q�,�kî �{ be�/1�K4����{����"�r������X�U��x��$:L��+i;�,^L�g��`�Yp6�)��cr3TX���Yh���0K�(Ȼ�)ODQ`�A�<�����:������wDD֘���M֧ֆٚ��Je���_�U��h[��e.=������:��a�(�,hr�#�gِx����x�c�MG̈��ML RM=��h��^����N�	��l��@�I-%!�y >���U��'GC��*��#�`��9�Tk�#������"����=q<�)�S�@�8��X��&2m>�j����t[�	y��E���8�KtBMYk��7kJ�|_����!��Џ?CK�/�%E��W�Ά�����C}�+��F'4MuU�\�;
�6��c͉+Y����,u�� �����@�ո��S&��E���� q�}��M���R6d� qD4��:@oa�ם���,	�����6�l�_��u�jBH�����H �ν"�E1n/��8h'������_�cS�ڍ�Pg��jO����@� H��;r�Z��ɤE�����o�r�_1{��'��J�}4�;�O����ČmG*��\��]ʯ�sY}X�څ��R4����j7�ЬI������s,�	f��&���|X1lf�6�=o�ˌRd1�9�8�]�h��R�X#��5`Ev�TId���ɻF�4��d��h��wM�O.��s�>���8E�L�jK?Y.u�c�or9���gOX:�ȣD���]n���hJ�2	��oDiW+:�央��@H�C
,���|�]����{��Nú��'�R� /�ZŘ�ɠ�8��T�i�����[�G��z�0�K����|U��ȼlr��Z��w��A�;�������-~���w9�h�R�|���/	�DB	���B�:�Pe	�0[ �c&��	h�l	������t����%K��~1݉������C����АD��p崾?]��g<�Bw��4���C�X�����[y��@ڢkˡ �V�cv#�2n���V������3����ǣf+���Z߈;ʍ2?���|`�C�%>��ʬ��n�I��������$2A
ަW淮��_0I3O�#"��3�]�7���3Ƀ�^�1�;�5τ����<��l��10�##I����}�!R�oG�Ρ`�{ǲ�1??�۪{����<5Ȃ�on���eq�Om�)ʨ����L����8�u�+\�H��~۽ �b�6Qh@�	��{���FGW��y�Ѽ��I#�&���������K׸�\��
��lD]��Y��*n#Ú�L{�� rlL���������&o���=!�w���y�|����\,2����&��W��=�=��0nA��ːs����Sq0��9��|�_����������_�Hu� e^��~�G����Gx"�w�]�t` n�L����s9CY�������8y)���|9��Ұ��?Q��r׶��'��Żs$���/�=�:#�S��9)y�/��e��2�[h�ȍ�DB_&�tpeɻjB���c]w�*�ς�~LD��/���S����m�K�^4��7D�2���M���f�y�)sF�-(;w�6�����`�ڜ!���i�`]�Ջ�4!&|��y4m�
S]e�1��b�؀�O�xX�� j����9����<1��F3�����"���I��ݺ?*���@0
�/��8*��(�H*Wv�6v���S �g��l;��I�:�MC�L,���s��%����P�r��dTe(�O���4��->��6��G;>��W���*�mՀ����@o �8���P]�]	񶘲]�{�*(}�ȗ�{_�)�*j�U��_$��;���R�h�U�N*ɸO]�(����[l�9.���� 7����&����+�y
-�yv�܅�l�''�i�Lf�ѕ���B��X�Dn���:mkkB��8=Nk�j��c���,�$�Y�����NyZ�W��t���r�Q����	�r##w�
@�X�J��X�疖�^�d���/����D��E�UH{I��Z�Aw�|�5.�������5n�<���EJ�|,����@�iL���oU��Q����)�>��ĥm���Rd501l�yI��ɜo}v'!��%پ.k��k�����C�33f�ǻ#�'K3)M�ViMnP��0vX�[�	=����3��z8�z.eq8�%�W�l���"</�.��f2\��p!��z��F��n��[�����J����a��D�x�B�Ш.�3����:jU��!є.���Z�t:�]{���)�(�-$s5 3�'I����nG<��H$M*2���G����efƹ��U��h2/?�dv)�9�0{K�_T���$��*n���K�i�K�qiix]���	(De�K����Nh��Cͦ<uHѵA�ޟ�Bj�����LŸ@s�����'��nԯ�8�e]q�v!p2�I��I4��PP8�7���W�ݐ���W|��o��.:���%]x��Vȳ�'����X�I��a��.Kh*�j|�v��zm~n�f� ��{[U19�\$��<�D�%�({R�:prB�!e�1J�9ض���p��i��f�K��$��_��!1�`d/�q)k�8; �����W#�K$����k��G�=f���q�Ԗ�i�[�&�	�t�0Y��_�j����){���1}ͫ�	�զO��?�F�J^��ș���&��贓��v	�5��
K�=g��<�g�W�\~�,��5��L	QH�3��t�ke�%�Sc�5!5�Ν�zx�15�#%l=^��B�E2G��H�7񙱯��#�L����J�(���NQ)ן%�z�<�0!g��^S��֖���ږ�	C��Q�yxpz�@4$���{�l�����ѸtG�oA�.��:� ov�-=c �o�>���W)3Z�s�0�A��2O�l˲���7� �#3J(�D;@.�6�﷦���$|��%���� P�vdJUu�+�bY��Ȓ�H�D���p��ʢ,XX�5J��Z�z���?�u�I��ĕ��ۊ$G�m"
��u5a�<M�ctE>u}qK�6w}�m�s�o1�������7�_�r�vp^��C�����j����-&h�Y�Q�I@[�dB�G��M��u����t����o6�$9��]��Di�2�f�G��eәn��$����*�'����_�a�w~�[4�������?vI���4�"8���N}���?C���j5�o�X��M�,*�W�/��^T���w _s<X�S[�̲n{���YAB��W����n�Cf�\.�����f����V�k��_lbM�jaŝՈ�4݇L��k��+�zX�K!o��{���#�b#^zi��w��d�f�n�4Aߛnn�0��h-��0������z��;X,����G��AV~o��s�p��Mqe����mx�v��j��d$��U���$�Hv�OE.�+ o���8�Fl3���m&9�mb�R��<u'�s�䄎��?L�Y��G��#ZX����{r�]�a,ʱ�A�(� vG.:�Q{H�3�l�M��
�s4
W��7��LӉ$�F����S4�N}@՚�6�yO�K���B�>0�0b�i�:6�"�sIV�J�h��|흸C��t�+�N�7#���E+��v�"Mm�o��5t��cbH��:p�aX lv�	���������c��~����cE���L�-�R��N�]L6�d7��:��ʚ�0}:Z�:�%��M���O�k�<����~jl_�� �G�&Ln�����{h*�*�|��hIK�࡟-�W��So�h�o���d�܀CUgY:{��l�Y��n<i+9��0��Rsh�esx��������0���p���[nw���m���mAT���Tӷ�%=L؅^iҢ)�*�_)mV!E��7�&Y;�l���Y�^ ���D+99C��)st�q�'� u�x�U�)�	s�0����7�2,���L���c�����;��=b(4 �/ߑ��S�9�^��������m���\��kF����U�|�,D�8�6c���#K�WX*|oލ
v�P�m2�N�#Ȅ�3;�T-?J$���τf���	������ ڴ�e|�Kg���9��)I�"[;\�U��iW@�)3��� ����i{��02�cV��E[�.���T5�&�yˬ�t���mQ�.Ŧ�]��zMLԈ��lS��>v�ܪ�� ��Vٜ"_�K��aӫ<�ħ�s&d!�
0�t*U3|t�ez=��>�4�&�9��66�:Ϛ��I�z��$l�l��א����P]��8�W�z
�f������ҩ�P�N��΢ �rU4M�f/A��wi.�����ОTҍ`� ��С�6�#1�iۑ�Exㅘ6	��w�A�~H?5��zvY���r)��K�Wy����ٗ3ej$U�x"�����J�L��y��^�g�g��/�'��^�א��s��E��9Ǘ��ꗒ���I<FAu�\A܎���0�FRL�Z�`|��e�@�}��~D����8o��B+,,�	�P!�3��.�WS�oVʣ�g8H}��L�ةn��@bas�����v�'����.L�c���)Ȫ+�Q�~h�m��\��|�~�_i��v���.76����w0��{g��۵T�7��7���b����V�戯Qw�~�ي�[�Tx�_�s�t��8��5���S�s3TP6����.݉}�Ye?�x�^A��ճ�~�kM�,?��V�i��H5��s�F�j�}j��7aBR�#�� �`�(=Cf����E�Kb D�j��R#�犖��fT �g�+E�������qթ׭yǾ��u���d�v,��u��V�X[�*�u��_��3�V���w��|� &c�VZ깜��r>����������WԚ��Ө��m�z.��n}��-�׼�������F��b��Ң0��U�0�x���x^zPMQ̖L�qjl��|%��ٳa`_#+��Ib��t0�$��WB�����&K�8@��Ж��ʵ�R9y�WɆ+�����,�'��Φ����&a�ȣ�CB�1�@�ť�<��kP�Wz`�>>�Jt��9��*Р��rvwb������s�4��O��	�8ϒ0�Rzi�ԩ��$�R&�HRS�*�E���)8�p��3�/�1��7������{9)�y�~g��L�YׇR�����%�0y	��E����?_���c0Ѕ�˿�?|cc��i�iw��P0�ˑ����[�9U�Fݟ��v9)�]i���h�hW��-B�&�L�%F�4��P� JF)y�*h�/0ܴ�L+��x����Z�a4�ꗝ|KZ.�={�XS��^�yN������8�ʵ�XC��.�Z�����~a_��ډ���x�+��;����h,������dBk؇t���?P��*�J9;7�]�^��Z�<w�{�m��ߍ<�?�y�8��R_���5��R/��$�K��@�/v�h+H����x��f�ú&l +�Ƙ��T�'�������~�;����=�O�E)�A9�/U.̬��U�4���Ӽ�W�_ŀ�d �V'�Н�u k�"Un�����3���"��ڛ�h^��W�t���ͅ���P��8��}]?*ȎY�p��y��-U�VX����x	�0�'�]�� b��:Η��{Z��͘6K���ǉ��s�܀��@����hWϺJ��wخ�oB˷���F��w�)�r�F�H:O���Ǘ�!��@�����jÕ ������ 5�J�����`�(1�W��_&����Wc� �5Ê�Y�9��<~�Ս������pG[�99hH������'k���0ldE���p�W�p5�~pR\+R��R���!�k.�S��3p٥������u���Z?��Dmk�#�	Q����F!���X=P����ė׭w]��o��NRl��}�}|�k�oTl�	�Q�o��hET�����s��\���2X�����R���f�d���R���I���NF������c�n(3N*�Bՠ���[hmfEYGI;蓓_�f�<��b���&&��료��E@Kc3��F�i�EP4�tN����JP����k�O���zJ�V����4	�ܧ����1��֐�]Cձ�ڄz����F��_G�5��R9��t2G�i��4/�	"��n[��!6��@���ip�GdL��Yn,m
�:ä���g|�g�U�,7f��S?��*��)�m��o�Z�����&W�4c�^о��������֍e'���ѥ������jr�O������Y)w*"�P �RFi$n���;g`��r~�Md��^|(0�&���J%hZ3��a�bs?��c�k摃4�:g��;!�H�J���bh2+Z���J��>�X�~59�4�B���x\hi�Q�¢�_;3$�`J�/-��ϊh=�ޫ΃y���ړ'��+Cm�4��]d�.��`f�%��B�\���N�q��7hҗ�ǋ�S���������-:(
�b�jp,�_��?'�yT]3j��^��nͶ�1zWI`���������7���U7}�׶���a'�M�a� ��1���P�T�zeHB]��ۖj�C�+?+�rtI���DQ��g�$�ȥ`ѥr�����#�i���|�{j����"��$��\L��1�X ã����y����j ���L�X/��Jv���'���b��� EhR9�a�hd)p\���-Sy7��\â`�M�z�
��!����Xħ��s
:��2pD�s��+m��P��y��^g)��<�a�QIK�OZ���JwѡZ�}�fC#�wf����I��ۣ.�9�q�(�>=)���WZ���)d�ƕ.H����
Έ	������Ϝ3�ND~Cf����hћ�o�H ;T�!y&�̡���O�{��6/b�@���vwx��@"ܬ5m�.�OO����*�6��JZ�@[�l�XP����j�(��?-����=/�a���|��0�2{7g�c�V��[��|%xc�P�U����&݄F�
�fT�90�{hn�945g�$''���A��c>�}[�W���f��� ���Xh�W\B���q��*)� (�����\����!�J��!��*~�5�RP���l�W���-��<��ta�)�f�fA�v��?H,�s�~��!�C�4z�o������}O��v�lG�-j�����`�oe>�|�Z�'�wS፵^���KL����nW��n�[�c�/�C��?�����^�7�O��ˬ�Zt�ښ��0�+ba� jֻ
�?p�;L��1pj�$#'h���,@Myڐ��V����*��YN�
 �c�6�`L�ۅ��T�(�)���Vڏ
&��%vxYv>�;^�"��exo�)�x��)*�5@�.�^��c����wsS�\�q��@`=씟@��b�5j�d��kG�85��o9G�2�O ���rI���������0	�K�Q-dvK� �~ĳ�A���	,�g?h�H������ߦ��Yl������Fy�շ�)GCLu¨�>�PK�sY����2!�I�~�:����i�����H����_f��3o��A���Jj7��AƮ��dY׏����u�dK�	�(~�t�)B��}(ʲ��uk�<�y�D�{����Ko����'N�������U���*tIؘ�-?�s��Hl�G�;s��Ay����qy���#K�js�+����u,��oOS(I�P:N�4t	/P�J�r�����L��e�C3ߣ��g�����}��IuZ���Mi��PC�ݢ���2��-)�ܯ�1C5F�&H�&��x�# ��Qe=�
3]�i����̼tKڨcOk�܋p#����I�.�F�<ũ�����o���B���א�'��ȱY�.�msk].��E3*AI$Z�k~��I��r^��U��uY��7�L�.q�4��z�0�#2������/�'��	��Al�?ע�Ұ��^g�)#�,�y*����$�Q��qjþ�d��H+�Ah��&;�VK����Wd�	0�L^���0J�w�C#�L��В�I+�A��	{��bb�C���X?��Ҏ
Z�����o��lz=
�o����)4��;��e[vx؊ñĩ�tR��m�n��&*�]�ߒ��H����I�kȫѺ�����{-:���C�_��Z3�o�:dS��#Lk��=Z�0�<���\��.�7��hT٤tÝ�Z��K���aM0O�p�����ŵ1��I�+Rn���!�Ƽ�llDS����Ͽ��}�2��d�gҸS�єR�g�`*���[�hq#��,���ڀ;�VX�iX�R��/��Q>y��.��;�¨3:�������T��j����wŴ��`�G϶�}D���:�=�5��'��P�����g<��}c�����\E�B˲�%�+�%o��yS-����c(����>ʆ:���6N�By��33:����y�D�IX��-������tH�͘��pVL�\�@��b˳5���*yd��{r�����EZi~��L(�Y�J����K��=��҃�Yb�;S�+�,+�K�a���RR�s�Чנ�扑t��:�Ƚg�_H[Ͽ��y�s�K�uB�
��{�kH&�ߙ��G��v^9��듛<?3�����06� r@5���]���-˓��L$�TU� �3�b��+/���n���)���'1���fb]�Z�@=A���W^҆���Q�P��P��u����	��FYQ�����kH~�;N�5�ŇΆ�`��s��:��p�8N��ȧl�	D�"	�
Q\$\[U�X��>�D����sR.>��g9�47� �������T�"�ߤ��cs�$����N��
�'qX/������R> P�Y�6ř��\�`/����w:��,��H�8�5�	[+̑��ZP9]��R憨��A���".�;Hq�iMd�*~|�eO�S��pm�:�&�`_�'�{���q� �#�������k;	̶��߆�ЕI��-��9\*�@�|G"NvtvM����ȥ(�����%QcYd���y��{��6than Tӎ�d��|5��@�%�iP� '����:�"�\��մ`�?���H�ag�����Z7��6Ԛ��5<!�_I4���[1��6����b��m���o�?�[�E�f?�q���5>a���ִ��9̓q�;J}����.�R�9\Z�����BNSA�c�?7~{AF8܊���P������'3"7%��t.�� X�fYJ��0!C�z���c;��j�Lq��j3弰�.�4�F����٩\Bw�u�����,mrW|\��P4���X�N	��}#�:
� x����HM��D��9Z
��{O��"N�-z�(����֛L{��I�.�⫆g���?�	�xݦ5�f����Cx�a�����s���q,i?�J`���\��򎞅�:�ӏm�]�<Uxv�s@�q�+cgGE��*�������Ȱm���+k��$�썋�7�)i��� �t�g �:Gp����u�Sj@t�?��K_'%O6x������a�E�>)h=����t�J"!�!:�In�Q�T��[�Qo7.���(�I�yXZ�Gm�����6�U(�4eW�;��f�t;�EK��~h��hP|ᄅkdO��}�uweC�Y �"�2���?� �n��/�"��z�瀰����#���*��[�0�u2*_�Vt�QQY��]Yh0�o��'@�L%�I��CYU���n���n�Ny+ӕ:b��9f�&��-F�z���V<����\�6����'�Θ�X�V���.!6!�#���oc��h��u���cC�$���]�_�����U�w���f<�JX��n,�]�!�����[��~�6�dc -��C��%LNT蛕@�`0��!Y\1
