��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0[0���.7��9�UU6�?�M&A�1,�q*q�	:���ъ�%��*�P�C�Ԍv4Ǫ�����O��s`���w�9I�-ĳ9��*��y7�E+��!pCa���C�0�D��j�cw��'!�6��w�ƫ������d�I���Ν�~�9FH%	����i��k��eή=9̎v>q���HҎ�#�#䝭�Y{�N����C/G
��lH&d�9	C�ɂ�C��vʍ�.�����2.�K�'x�([�5�D*��F��CP�Ǯ�{/��������&P��F�ښ�>7*%�5���c�Dt�pa���q��&E� aN��}��Н���.^d����|!��a+fc���<gU�co_Nn����T��ؿO6�/q|����_�F�S˪}a��:o��)}��v����E!�"��͋S��8�����;9�Gӈ%�ڶ�Dq��]���2���_�h3�90_z�!�"tDq�)&%�飠2�i�w�{�p��qnh�=}��	�~ �S�2U��[�:L��+��XJ��y9����?P3{��UF�
�����zU�o�*bʢ�F�(��@r(���<�D�b}�v�N/��ͦ0�F����+,6�/9��$å<���(�"6��ۑށ�� �\{�JF/�{���yC>��d�.?�������$��/^>��Mn�O�����0�j���pק�h�ڴw�ӯ����Y�z,�J�p�`n���j����i�16@��-����<����1y�J w� �xo�'-G�1���{䨹a��0#��k[F�S�v�A�oaYF�u�/�*Õ�̊� Rv�h4����G��Z���9U�+��h3�@�E�������pk"���:2��_M�6�2�S�y���Qݐ��3�13�^IIE���p����~L|���!��0;�c�L�yb{�wF���9T��\�*G����b�g�
 W/T@f3�uw���ۄ��mj��6�&�����	�a�Un&SUn}�hLf���:ܤ?u��tG�4�4�%�.댜�\���v�է�W�����v:�M5�V����H>-V'�w���ɐ�0)h�H"*�&�Z�Q�퀰6�q��� A��Ws�C,x�i\�����+д!l9I@�ߴH�Q?����y���m��(H�q�r(�h�fݶ��\^�R|���	��q�#2B������*o����ٕ�+�fM��^i0��ң[V{�#4���M��1���)�@ٚe:��V\Y�#Юm�e�P��F"S���A�*�f�����)���s��E+�~�9]pܖHNs��� ��q{�>y�B*�b&huD	ؠ0>N~����PΈD�{tծ�]�L��	����|W*�/����v9����p�c��)��d�-����na�����>b�ɧ*{')����_+�9���P�zE2�H���e*�hᅨl̓�%bR�
R��|��
���R�b�rq9�x�����`z��)ٰ�6ܬƌ�G/��B�},8	,�&�; kJ�=.��K��F�|ۛ)tq�^��7L�[�Z�LS<����Y�4a4,�5�yVK���ס�ہ|>���B���?I��cZg�i�V��V�J�-�~ ���Z�m�bt;��b&��S�VFWi�����f#tG��Ϡ�+Xj�-vw
�< ��r��i^{8P�GP��V�g{I+����tlc\_��\㻒] S��V�$�(�5Z��ly��B�]����4�����|�}�B�Q1�]]X��n�DLOZD9�A/��KNpbP�ς�E�+q�y���p��~+�<������@FC��Fɡ�@�z9���x�F�� '��R���o/ic�gB�K0d�:Р*�.xB8pf��y �u��(#rud���Zi�'b3g~��uhɣ��G֊/,��i��'���eb����)��@�6|��;G)�&�%�O0<�U�d���4�r1�$��T\���6�0#N����ѥ^�bQ�G3�Ds,�%5e�5�4t�ALG�}6����S��2�SJ*�Nw��e��x�j��Ǵ�Ǐ뛎�ER�$����C��ȃ3����	=�����t�y�rrR&��tJ��*q��l�=�M�;b�.Y��
��?F��I��}�\�&�Y$��C2(�ME���(g=��L�v���������G���K��a��J�*;~J(#��l>f�E�O6}CRZ?�$1��?A\��g67C0@�v9�؆_C�V�u9���TȊǙIh��/����n�])��*1�\�����`����F6ɦ�I8M�cmB^���#a�0����V�-�!�a��������DT�q��0�Dl0��w�%� V������i:�3���M�8���q!�A=�Wj@; t�~h/����ߑY0�� aF��L�����ȫRZl�5ɤ�)�'�T�^�r�8�N���$XxTe��Rx�p��Vi/��I�)]>�7f;�Ƨ����w<%3��	���!�o�%t�x��6����D@��]B:)B�(o�iy�)I6��m~�����!�e����|������A�!y4'�J��0ݎX�N�:���e��1�����4;��mؠ���I7M>6�-U�k��["�u������* :����kA�&HL� G\�=7�85�9�ج{"A儤��8�X��[m"`�Q�4c��.\	cr��N3�a�HG��
��a�W�ڴL[������X�*։P��_i?}�/ִ~�N���j�3�S�#�Ǚ�d�% 3��L�X]�'�2�T�!���@���q:�	�j���ft��m��b,*���f;�DmBk%8?�8�-uÆ�r�X�TN��Tm����Cr�Zi�w��8[���`G�5Иo�b�\lj�9�>M�D4����ٯ�P���ztn^�>p���B�OT�1?�O��9�X>J6w��K����kW��K�UMQ����:L��Gl���b��վ0���Z��
Ȯ.�o�:%s?]p��H�B�� +�~Qo�أ�	��簊�4��%�����%�o{W�k������q	(���`�;��\�8�,�6�9���'R(���-q5e~�@����s�Nz� �U�m�ypG�0s�Ye�D�N�
Gݑ4�M���^�|��@��Y�Hl�+BX�nsl��߽�
��}@;,DH0�#�*)�%,[�X��'c��qS��XΥ�&��ի����@��+_E:�gWX�=�]ܯ���րç�Z*�!JY8�ef�b.:���2�M�w[J��6���,|�AUE�lmr��(0U�]����z��yJ��Ʊ/"�ߴY��u+En�]�+d�����*�EeRT�*��xA����%���c݄ʚ���S���s�vh��#���xB�9��q.��pP��tS�v��1�$z�D����Oa��2Ծ���A��یkoT������N�)���כ�>��=!OS��gm�p�Ӽ�<��8�i(�T.o)n��Jj�'Vn��G�����{�i+P�&NVFTP(����B�D������O����{1V���rx�MR\3E�ߣ#�%�D���]eX���|�e��j���D��~���g�s{ن��4���3����i_.�-5C�6M��3�R�wjQ�����&~x�'L���X	����wd��9��H�e��F��ƞ�ʰ�uY��m�lEAP4c֮L �i8'�{y4$K���Ԏ�;�c[�:�w�.�ѓ{/Nv�!������>�#w�Wj?k#Ejֵ�J��^ �I�1�<8��\fdN-��Hе1�'_��
=�:�/���"�Ђt9C��b�n҃�E���b3�H�wb��]V\6���:���(\|ƣ&msLA�E'T�E=�}�T�wWo�v��H�|�_����E�����_�
�[�S\�G�i������J�:	��C�Lk«���
���Iw��i�OI��%�JcփN\�=�>�L�n���8=`��j!E�#��'[�wQ�xS籛[��bC�E��AÚw8�|\��s
��>�F�zeD�8�j���[Jk��L��{�B�������Db��WTӳ�M�������~��Ɵ���^/l�"[���v����\{L�&��Ԡ��c��L���Y^����6Q�kL��r8g���uω��K��K6V<���KQ�Թ���K~����b⤼����[�J	Ђ� �S?���>��Qveb�Q�bù��C�9�2Y��s&�P�(�V9�d�)�4��=�S�A�~���.��`�g�V���+4��q��iQ��]ɺs�3�<���9n �y<xn�PL%0��k�]�D�3��R���~��+��TD[�a��s�C��'�iu�X���!����K�� h��Bg�.�;�k�@vN�Y+}'i�V�abYGq(&r��{���ߏg��v?�xě�ݷY�z���%Te��f���:�N�@x�Fu��8w�6�`�&�w���&�d)fBID�kqR����5R�|�d�ܫf��ꨕ��q��T9v-�=�jf2���~{X��喳�T
1	��1�vq<���}�u��oP�Ap���?k1����|�t��+���%�����j�$�.�	�u� �X�t�&+���9��K|GY�X��D\���}����L�)��
�y.]�ZՀ���K�Acљ�����-�HL���q�Cz�������8�A����PΨx<�RVJ��^��Aa�rX�n\�?[�A��V�x�j[1�Hi��),��?'�c�]���i��N�jҗ��������8���}�$��߉Y��x.~�"9�����rֵ;P[K����O��m���sp�.'2e���Ĵ���O8x��ŧ��)u Z���o�_�=I�<���!!H8'��.���� �t�����W���u�>T?2)�� �v�7h���˕7��0;Ȓ������ս-���E'��U��9���Lg�;/�ߑ��Fٵ�P3FC�XJ��w�6d����(]7�-k�G״_·�5J����ެ�t�e=)a
��p���c;�X'&X�	�vd`م=�i
02鳺������t�j����TĤM�����.�R�$�Y���Ts�t^mt=���"~��#���F�v �܃�h�`y�_���0����hK��ey�0j f~I�.F�B2b�4��̿���X[��ʥ�ALx�ڮ����|��d�`Ec"B���t:�|�{���#Pߑ�,j��
��|�Pj>0\���P��ij��0h�ɧU�@��r?�Ԕ�ݍ������{<�Ů�:����1�[�nB��:��\9���"]gk�%����R!�JƇ�H�Q0���N}S��U�^��Ed{���p�[�"+��/0A_B�7������b�� �C�R��^��y�'�г���$�g|~��/�9U�T���@%�}!Un�C� %���q:�U��莬X�.9��>����Q�"}�^Z�q��C|e��1;b�=�YU��A-��W��:�1�h[_�ګ�պ�+�aY��>�Y�q�O�
��OP�H"�=�<�x1<fzsȦhz!���Ti=ćM�Oa�D'9�y�������r]�Yu�5!B�~�>@��Y�YYÖ����sЗ��9�g��s?�sv���{�;�U;�Y��R�1�*� �;��s�q�ڛj�%�˄�����?$�W�njR����0e%_p��tE�Fq.����O��ںi�C��Nx�0-,T$�T�_�	��,h1�}��!�� �8���t�L�A�Nv���U?��B:k�ռ�9d���{�d�?y��7�z{!f�WME-��	{b�]>��n_}��[|�7��)T��:t!��_cŒ�����1[LƫK�_�V!䙵T�i�_Y0M�{P}����;Q�����nݝ�/�Z�mS���~�]�B�kx]�c�0�"�>�Zɼ=��;?��L���Z�1�d9�HLھhJ�>�k�Jn!R�.��&6*GW�	���{#�|��qL��Ͻ��8�.�����K��3���x���e������fS����V��KK�?���Y��10�v���`�H S�4h5��_�DC|~!���r(L�)��(���1��O�R���t��;$�r��/@�\��4��w6`�A;�P���!�U��&xS�8R�@K�z'���62-��n�����pq>ȶ.Q]�Zx���:I��h]�%��*��t�σ�EU�A<U��?}���u��bmhe�Q2��QдDW6mE
Z;�fd�����g�{�U���-�OA��rg)qњT2Z��،���4_ҫc��[�]3�)[��<�`�ƍC8B��B�Jq��(�3�IF��X�����]H#�A|�Q~uY� 2�&D��$���1c�� U$�U��v��~�0�!�8�j55��:UP����>��ɧ��{�i[S�- ⼦�/��
��gZ�����I������7�n���`)8g��T����j�������Ħi����������c�%2��{�=��j��F:}۟+fd���}u��rvm��1���RL���#�%{F�Iya�u%Z[t:H�	s8_]?>��Ґ�V�-ݢ���@�]jZ?-��;T�ll�EA�I�t%#�B���˯��L��#���~�?|�|����>�����H�vIC�f�k��X�t�#x�1"x��Ў��VX�ve�7�����7�^P�s<5Fc�R��q/������i1�9P1*�a�����M��Zd��*~s��,N��W��֑�����GZ-�:^�	U�M�I5I��d��fN�wG��#M��3��r����c~���#.��Ҫ�Z���<�g�%����ڀ���P��k�M�r��T f�1����ׯ�RB0�Ʈe�hIɱ5Z�nKl R�],+J�rT�ˏmX%m��6V��+�lR���w��4*w��ĴT�{����A�[	d�Z��zR�M8��{cÛ�I��w0�,Ur�V���r麊�{�D�i�l�	��'�1ݫ0��k���}\b�`\�H����;��=/P��Γ��{Y:�HZʽ�5IW�2��ٹ��n�7�{���i~:�ۄB �k�k�G��J����t�G�z;��(�ַ��Ѓ�결(��
�+��pe�a2�ETƿD}�ٻ7��ȍb!�d�w#:�Η |������|�tI��Á	k��h��Q��a70nє+i�EY�ԓg2�	��B�\��L���"�x'�d�K.7Pfd�Q��_�`m�jC�(43d�CLraY��s�z�Hv4,������?�8��KM�ƹ�%�~#�����fz������:Υ�(nӰ�ɮ�h�Ԧ�mb�q�,�6�2	f�Njp��4�f5�WIy�e���I�X9�P��g��JNw���2�Aߍ���%��Z��WL��ш��D��{�Ab��1��!�*��2h�	>իMG�n��]ZN=;�b2Sh� ��HP�~q)$�t�#T~�v�޷B����N��� ��a`�1x[�9�B�!��"�K\�d�S�6�.7ЋJA���JP~KO���N¥/�ft_6ǓG�,,|�����C*��1���{�m^|4��X�r�yw�N][+z�j�8�q��D�C;�زƱ�|��Œڞ�YfB����Q��E~�pyG��Ӂ���$��1�rD_�d�ך!!Q`�'%�a�f>��G�Z�k�M?�4CS��Ӥl���6z=�
�`��1��Զ����[]���6����X�k�҅�z�+���8�é'�q�5TS��U�a���z�dC��J������l숆9s�V�@
%
��4��%�7�u ���iu	`>�E0�ɤ|f_�S���aL�^��E��L=�����h�d��F����2��h�d9$�U�fA�l�\"MBiЉ���:rK#,�R��Tt���\Nt,|U��^���\t���]�Ggn-�{<�{$^���+�W�΄oY1s��:���!
���J����Ե8���E��v��L�괾�0 ���8EJ7��vy�����*����ԏAh㇚�^TY��<n�@���+=�kgJlZGd.+.嘇q��$[���v2XBTp�J��.��5�F�����P���el�>r��[o,2&Sɹ?��TrQ�����y͌'+R��r�"����G	��A{h�P>c��@#촞S����	I'/����a6>�`]��֍��Y�ڧ̫cֶ� �_tT�,O��&��V?F��#Z�?1��XR��6w�91���[b�!F�'��Z�3�+�������q��,q:@I�.Ԋ(���[���G���aOPgߤ����;�^l�4F�иB6<mO��� S���_�{�L��ZC�t��{�߯ݍ��#\���E�_��I��a ���XYN���S&�jѨ��B�P�iFԔ�l��z6�`	���O^99���j�lPq��q!��2P�lS�W��82����������u���E=���ZfF��E�[���Ay,�v�
�� QPT���bZ^�.�*� �Q`�@�,��0�����B?��z��^�,�/7�u���Uܻ��O�+�V֘i@�����N`��ّ�~��/tn�Y>���t� �D1�I	��`��t�f�j�@�����g��O^�q���f@8I�sv���q���GE��.��9���4�M�$�e�'&!��{Z�5���%d���;��'�j���̺1u����Fi]�=R�6p���P�MMB%9�e	��q!�Th"A�:��w����q�Z� >ٛ�R,�">�ғW�tg��ϥn~[�������v���O�{w�Ő9��=�[�sAT�7���"���������u��W�w��n��s����Y�E�6���A>��d�{F�{P���`�e��z=�����)�}�Z[�8â�䛑��e�K0iOd��g�e�S�
�;�&�Y���Ȏ���l��u�<_��{q�Ul�ְCy�����3KޤZ��(v���S�|ʖya#پN���sЏ�I+9��k)^�b�5��y��G[/���h�3�ms�B�>��� �3����T��AcM��=.E�7���`]�>��0�s��"�HT��tjgtif���FU9����@��$\^d=�JB�	�7x8�t2.�����a��X�&���LS�G��� �z�Q�.NZ`��4 �`��°�1�"���i��`�dփ|�Qg��$� %%�JN)�+�4����E�H�����&j&Al��б�j��u1Ob�
 FNz��s�F����ɡmi�4�0vI-�p����3���/kO���O��u7?�m�a�[էʕ�11/V�����L^|�<�v�f����N��_�����eJ��^;��sw<e�j�����y]�x2�d����[�K�w*7Zr@�NK.��m`��
�)�?�����˫&c��w�a;�g��,�T�pPLsew3��#�5V!t��4=N8��I�9l���I������EO�=� 5��,�ƶ��G��$�� ål~��U�m9_�\��G9�a�����Y�8/��F��t2<����d�2R�U�*��(@��u�$/���X �l«Y+qgN8�$�Ǎ
'pS��mCJՌ5��L9��� 3�#�r7t�d`;���]ؾ2M}�-s�雈+9��6��X2ͻ��HM�pK �D���Un�+����
