��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�Wo�x��s������Q4f �a;ON5�/��W�
��Ϲ�(���r�85�8{HcA�E�Ӑ�
��#9��:̍|$\�Z��L����iKT�dӞ7�02H��:�x���s��^m�Rq�y�}P��Y����3�3e���-\4ZHE;/ω�6}u5r�Yb���<�6��z��NG����pW�*:;l2ay�V�[�����>m�m��Sk�@�� �ͺ�h*��AF�D���"|�A�m9�a�"���:�#s�,����B��15�yo�J�����$s߼��
�F qY��yw�5���#j��V�cd���^z1�5�E�=W��6]d�k�;K�õ�Yh2�OV;P��,���k����V���
�s��^Z���F؂������ًA�Ȅ��iM3������)dVo�|�����(7�gѴ��d�r�]E�>�맑_v�2�F&�^b���	���;�8{9�>��Z�^���W|��h �R�(p9��g�j�_��j�ўn2ZO̹y�s�2�U��{*tLۡp��)����`���z/�g����gK�ƾ�꺞&���׿�;*���q뙐|.|���� m	��"p��{�A�)�죊t�!�{`x�!3R�:���\���đ�e����}��Q�?�v��)��CH0��j�9Ļ�����Y{f�d�պ�qe�S�>���߀'��a2�K싣+�ش�NQ������<�&K�vO�%G�Σ왹�@�"�B��8MG� �Q�6�=��,>�.�����g�� A�]�QȀ}����4!߶���G���}wѬͲ��L@�2�i��H�4멲�ɏh
B��޷@U�s���,�GU��Ge�
*�n��1�Wf�m<@w�ϵnW��$��sȧ����0;|�L�}��:�Rjk�=$ڠ��Eu�����˛�F�6F�&�$r�w��Lض�Udf����aSK��ϊM�}D�$�Q�^��z�Ҧ�5Ú�Mnp���T`�����Y������"�2"�VG�NRj��
�o��@���[�b x�ǃ,V�`�� �g��# �юm�Q��t&��kT���Ax�X�8�~��*=m)]2i�m��h��ͤ��朐��G��Ǒ*�� JN?�7��	ʹ�3�V"�(B�Ug���K�8gi���w�3��<A
-�*B��/��S��%ܫ���b���ܪ8�4x\�zd-ދQs��(��(�b�^�,0px6�|���)�< @THԨ�%����3����_��=C"�9����6$�b�e�p�x��#A����Ǧ��8�B-f��)��	�����p�h�
>�[J�K�UTo~�FV�7t������PXz&tL���X�?�0q+Ԗ�f硃���}.�S��,<��9S]E��R'vmd"���6B"�H�H2����L)�$�Vۓ����B5ç2]����j�߀�cyF�宛���:�{2*u��"b(œD)&�����?�"7�A�^C���2|�`�Ц�	��-�p��ݙ�j�^�$\�jX.w����}�l���"�t�!�YK�4Y"B���p�(�C�_�da����I�[��O�P���:Al�V�������*A�%w�#x�9�*�1��uR�hs&���m���͵��g�ݰE�]&�Fp�͢���Zؔ�p��W�-Iw�+E
_��h��P�,GU��0�����r?r���9{?cdp`E	am��aVRV��{2ǡ�%�]�ҷ��ߝA�uTSɥ�~[ u&^&�Xu��)����h`� ��I�{Q��{}�>;q$�a�xϻ)1�� �yzM�L�}Dd����,1�q�S �O�f�ċ��F�~�+%������e�EVp
��Kq�BU7�\��$��emNQ��h��A��!��������A�Z�''����[ɥ7_�uV�c�w���$�@O�?��v�G��@+�+z��u1��3��t*��08T���0�2g�E��[I���eYB7������f��SҢ��C+��A�����a�$\��<�������4��=F�]Cu�=��g�$�_)�1���vx::��z[u�(�Y���x�5� ��ۜ/������{�[vO0�c�,�?��iD��Rn�sGw6z�����ʸY�>q�	���l���ˢ��c��XI����
��qMVϫz��d��� @��S�Oj��~^y0�c����Hz��떟��p�:�U�&	S�*K�s��gp�X�Z�'_b9՛?�L����R��_x���Sܤ�����'wTB���E�+C��ll�9P�Bl��d�7��UŜ8cq�9�Y�~*�p�I��a^�� (\�#kN<�z(�G�h!w��t�BC�f�R�
u��)^���7r�~{Fj]�S#����]�+�f�	��g?H�$!`�7ĔR�uu��6�{��մܷLw��K���&h#G�NX[%F&vթ�~+����p�:���:�{3�w�2�c��b��u��~d��zMŦ�G��"�!��%��㣘��+����&v�P 8c��)'O�$u����Hn���^���ql�tx�y���������A��L���k�{�'�Π8v.����R��AB*��*��\ʸ���m^8S�:���EVb�#��	�La��'����d��x2��iK"	���i���n;�sp��n��Z�k�`B:��H/��ݣ	�\w�vm+aRZ��BC!��7���ĀZ���fh`Y_k��;���~ieu�j�Gek"+�nr�����S�z>Ϛ���Z�I�)�9���0��֖ܸ20�� ��E0?$"���wGbd�0���d������YKC��4�@&D����p�|{�˚�H�~������%�×I�  �?��u�ct�$�!͍8�[R	��_[�&O*s5�u�TE<��L0�q��FD��sD%��W}{A���d������
Y�R*+����j��j������C�E�r�0�j�Y���fc)iMI^L��ܤ�L_�����\���#[��"��2�}[+�A�������Sa�O��F����}�(
� �Ɨ��O�Z��4���Їj$g��?�o�/�?��X�]��jyG�zbN��I&��e��Ϫ��(5ZMh���y���c��k�	�޽H��ֻI���k���z2d�d����`�o����m�A��tmrw��Ļ��˼��ُ����VQi� � E����	�z��X	*�ܐ��߶/��R� p{�b1AŤT�s�,���
ll�~:Qߖ�gbd��T�Q&Cu��(�M�
sQ�>S ��ð�m��)��'���.�۳���7Z�pI:��_��ѫ��^��ĵF����&=垕'�����xv�_����?j����pE#�H�O���襖�{ф a`"F���	�V���O�M,��9�8y9�.��N����k�Gt��~ޞyP.gf�D�Z��㓁�j6Hj�Uk)�~����t!�2:#I��R6i��ڔN �2Ā����Z`�}���p����z��3��,�/�}w>��i%�8��CI/-`���N�P:/�QX\Q|U@ã�JѱR����a�z�W�����{����Q˝{�:u�Aj+�k sw�����õ���~�N�����@�2�ȷ�9f�b�h�Ao��f��9^Re�$n�_��߈t���~T��>��Y�c 3!Ԭ�����Y�^
���� �\����}'��i��|}���u�4��w:bA�E�F���2��b�*��2g�)���W� �	�r�pȺx��SS���ծ��� �b��yAz��8��=s�#�e�@��N�I-��`�^��z���M�����n��x�F��ܬ�$�4eE��%<BL���}J�}ʗ|��f����l�4$}��;(�r=@�?7f���Nɀ�.����͏�V����=~t�{3��m��W�pk�?܊'Hg3i���j3�;��X���"�F��۷�厜ڇd�C���dx� :+C�J�B���DX��_[�&��Y�<6�A넖�/?�ɘ��&��?(��޹��''LQ}׌�7���}���BT�U���l߂Y�쟋VT�y�U��E�m��� )TZ��>���ƚX�Th��M����^1齍?-+�*O���7e�B:%�ʘ+5)/�d�*�s/��t*)�-�Z�����|Ϗ�@�C-z�Q�ebx݃5ӣ�u���?q\�?7o>�����Ed����pgB�f�b���vu4�m��m�����ʡ|�X��6��a�Ɗ�-�U�g|�n�rv��4�]?��Þҷ&�%�����_���ЕC�d�;�����ѺQ�s˂z��ﯣ&��	��h��Ǩ4�RfX���4��	|��O�H�pkRE�@��l�As�c�V4�SU�ķ�H��A\�J�:q�xZ��c�"�Ԃ��2*D���/:avj�૯�ٟ��{��g�Q��| 孛5�ɪ�ޱq3��p%� Z~����\¯��;o	��x�2+q����"-��?7�'�:��z�����J�G���O�ų���ƎoA�֬yĔ"O7R��V�u�-%�L!��cз�i�HE]J���#�X�c4D�36���<À5���Ji�1ᓠq�m�4��2�'����ҕ薄}�ĳ1k�B8z�_Q%�l�������J�o]����ƺ�F���pr|r3~w������uGX�JM+z�d�j�[�.���ظ��e~�:�ݭ���L
����JH���u�*�I��ɸ2�dn�w��"6(��������]�@�~I�P@���\���V���ض��lдg���g����4ORw��K�Ч�kȱ�I��~�T�����O��E?5�I����o@:��Ka�؏$�,�\�>7"ʡn��h�BW��٨%�23�"�%ɧs��W�������dk�P����Ƣ�����0,�5�l�4DD�u�E�\��z&�/v8;�qcu��-I�usz����3�MR�Fİ����Ŵ��3vB���n
�Э�)s .�^��ٗ;�P(��=���Ro ����~9`�aUڊ7{A����Mն-��,/�Ft�P'�a�$��ƣ�!c�tT�ڨ�r�N�O([��'��[��%��"�����k0T�p�21�Θ�@��U��$2�2vsW�W.&8�nǄ�ұf��~�(jz�~�
ݽ��W�G18��?��{n���=U�@q�9F�i��a={W�l��8P�$�d�w��!�=t�>r�u�����xHc���@�-ٰ~&c v������uu�yz�.�'8�����ۉu����Q���N�͹���zT&�l�L��-5�O�����f����@��Ʌ��+HE���y~��[�7������96������~[4��{�-�@��k��c��_�	5v�����I��ōS�r���c��P_��9�j���n�{L�փ�D���0�)0O��)w���h��p�7i+f`� �|�Zp��2hT��6_a����Q���\�Y���`���0��������#�dJ�p�li�j?���(	��i�^t �L�еE����
奘2
�xRe�q���$S�͟����dne'ȑ8��E����/1`�&N��9�z�����Ϋ���{dk�Џ�&��Es�H�qy-[�P �r���������֩t��"��O�pN�Ż�`L�^�C6�]`_-3���!y�T.��\U�	�=����&���exa=*��~��Mfk��_�|����d��Ĩ1RK@p���k����:I�%�M�;�!���R�g!D�kg�Et=�6B�X1~5�� ��3P�jq�ѝ����p�-��v ����jq��e�d�`�6Y*��;o��z���X��0�;k~������b\n�@}�n0Ij1S ���ԧ�������<%��Mj�yr �w���{9-]w�Gl�BV!�wWu(�)$3�U
=x��:��љǊ�I^�W%~�u��q��y���P�~%ș��GL�bIØ�kő�c���Q�O���� ���Yd����uGo��O'�Ur�$���,�hA�����~>8?;ˉݢ��f���$�vM��u��=�Ľ���[��E�5��m �ueo��  6!����#<��S}��g�#i�L����/;�mAI%���CqY�!,x�?{�mEh�5x0���2�EU�k%j�7���ś�W�ly9�r��f�"�#	���D{?7&ln0��M���!����= �[��a4~0�j��k-�S��ĥ�D'��)�y}v�&��' G>��[��׺ʎ�8����Q�Ƕ�o>��c�D�I�t'<��do#a�smp�Y�n��9�Ytxw�aq3i�ҿ����v�ۘ����_ ����	 y��}��P!@ϑTG�i��/1�ƹ�F��nxI]Դހuz��>��_�h|�������E�1���j0e��۰��'
��~�}��?t�R��=Q��Ʊ�D iY�|x4��ﬞ<���z�Hn{i%+T�yx��8�je=ڝKU�����W��ͧ��v�8zY��C�no�O��o�͌�r�����@.
�i�1�F�A�ot��3x�Pm�,�a��9�g!���ȳ��gF�aJ]����סq��Tc���>�%q�y!2Kz&�L|Ҹ��ٕ�j'�����[v�b�Y�[��xC\�@Ygʸ�.��
� 8�"#} �	Z�¼����y��Ѓ���ÙO��҂[��w�z�;�LZF�
�4���Rb��BS�X©u`烽��ن�e�=Я��̣��tul�T��s��vRcT�C����%�/��č��׼`��F�5�CUW&擆8�� �A^�]��-�q�|1�I��_u�T�,��<"1b��� �y?� �N�N�<����9ğ]�]#��s{>�.��f1�I�ujɢ���S�/�~��nٺC�1���9����M�4�U/�+�ɍ�f��Qrݹ���'���Q�<i[��3�5I���:
���B���z��]s:o�<���s�P�D,_�s�Ԩ��AOjTZS�U�9��ZY�G��� !Z��3#�?�w#4.�Vm ��W�~kߨ�\xJd�>{RH��sw�
}�FXO��[}?���	��a�����~	|�R�=˼8|[��S��q��L~��aP����g�uސ�AhN��q����;�$�}.�ie�Y��G�a�������)�v��5ޓ�gτ�_�Ñ�-���}3�}ɦƹrV�h�]P��b�8C�O��Ήӏ:���ܕ���?ژ��q�s�R1V���)�r��_ʬ�5,��~��b�:�xsE���7OE���\-i���N�܍������S=�d�_��r�&��
�R��F�Ir֡Y]�ǅd�6���K�(�ͥV-e
?����,���K8� ���Y�5�h��~�[`M:NC�����H6��2��ӫYU�˽�7���wܯ�%i%��+>��)�S��p�$L,վ�)"�0�C�a�~�mZ��+d>X!���&$\�WAr�Ц��=�H��]y
��c�}[��pY�д��Kg��j�����_#u��/�n�\��f{vc.h<G�OEI�3�����]�}ŕ����)�VEC���#��)>����&�p��1D�9���
�q �g^!w���gnС�mƧ��7�~�M��n���C������^�c{��8���ΐ�p`�&�����9հ��b�(]w�Z�;C���������BE~��4�����w�en]�v2�}�X�eP��s���]�����t�}�f��64h����vhoo/R���T��a27�'��U����,-������\Z�����w�̫����������Cqc�ҢJT)4��;ر�@m�;UG�	�Dy��'[ف�UoIȾd����+��cdOW ��,�\e�B�hD'^�������\��������OV�7=��2;��*K�+S�1oKw�n��g�	�;\[c���tĀ����Sv�������X{�֍��6��ҞCy�q���[h��,O�]��gJ�1��Q�xk?���< ��ݝp3B�2xA6��62��� �-�(X�k7���/A����i�,�m�C��S��"��{�2��G���߶n�1�Ʉ��8���j��H���-]c4�;=[Mk=+7Ch�s�����Q��op/ĥwV��G��]a�I��:�jd�-�	�=F(�� ?��S�ZP��и�LD��NL����JM���3M�����Z����_^��X��������>[��v�*�ӯ0y�})��*��Վ��5T��;�Xm��$(������1~�o|��M����v9 ��_���	�|U��.���z�;3�HM4S%s	xZ���]�0XH���O��S�����zB"9;i�c?�8�������7ƛ���/�_\\��a5Sh��H��s�V@��&C�4����q?�Ys$o�P�9��|�w�_�Ҏ��3%����D��;k�쩥m�>�
�����j
s�>��Y����bb�w|�f��+�� P"y�f�w���z����1��`
~q�Z������P�.~��BEg�(H{'8��E��豅0�?c��׌�tb#�uŎ�.����!^;K�(��q�L�
G酇�]�~��G|A�C�Z M�s�*��)���v��x;ZS��͉M)9�u�:yt�,�������R�?�G@L�$��-���}L�JG� y?�uzv�b�G^��D���[������@;;AL�1���f�� ��m ���A�"�L!����ٔ��BIj��1j�V&l�G.���E�-_�������ycvr�D��zC�$�C�B�0Xc~P[�8%��i�������|�d�lsn��E+r
�Z#1��x̋9�s���K���?m=��㣗��|Ȭ�l)F��^.�����	�Z�����!���L�?��#���0BͅP��HR�2���`����F�n�m67�;:^���O�`�9ɉ��a����Y"6,f7����$��%�X��GΜ����ߪ��= p�2��"�:C���U��i*�.�m�ȁO���H��ܙ��68���/��7QurwH����4���'�	vg(�#�V�2�x׵�S�D�LhSzԟ�G3����Ed��3����C_��~�I:)9"CE�g_�D�R��n��D�s"���RKU����z���HM��i��m:!u����0-���2�[I��7T_O�Q9v�r!�B
�����*mP9���,�ħ�C[��M��1��
]�v%�rvD������R����-ը������-�ECCh��Rjt���)�)i���=��,̓d�z/����C��R���E@�}����xps��a8���\��A��cb2�󠟔~X�c뒣�<�'�#����ރ��b7���a��ݾ{u}{�v� nt�_�Z� �ʘd�wpT=������p���R@�+#ncg2Ӽ/R�K[/a�X���&��ϓ-�8j[�Je,)}5��{�E���H�-n;M��7�����3M���ÝBr�-��ʂn3���#�K�?S��(��s��
�)ǏP�g/�{��K@<�d�*/������Ց�Ğ�a�-����J>)�3��K_�$�go�!"�h��H=Ǝft��I�d ������f�t6XČ',\�q�)Į@��EѡK��©�u���Z��T"+�����c��M}a�)=����zu���OV�hQZw脃��v�"�Kv��N�]$��o�ʈ�z%�!�@(�$_1O�!eVL��/C�>�~��qgf�[G9��}��,��(mX��x����@�r��~��<\����73��UWO��`��Y
�mR��qBh��"�� �vXaiV�.d�
�$g=>��W�F	��qO1iu6�xY����l���g����`�zЮ,�'7���b���!8S����f:R��������X����?���踈��Wp�5��D`�Y����g��b>�9#���B��<~� )����ȧ`j�w��抻ۏ�R��z�ur�;����p�Y�C{�LS����!��vS�f�M+۲�K��+�{ �CX;' 8��A�T3��	ގy� ��_��`�"S��a��Dw܄-4_<S�~jiή�(1����e1��0��޸P�9ۖ�����"*4��,���=?Q�h��{8�K;Y�K)��a.`�6k��qCI&>:�)�����ț-k� �&R�5_���`+�ہ�»9�A����_o�,1y^��1p����'��]���߽А�~x�u�jJ�]����6���`�6{A��_	Ϧ 5S.�
�������"�x �_�1�rX��l�����6�Zp���e��3qNl���]#�.��֌/��<� ��4�Rko���L����v]c�^m���nS?�А�z+�J"����?A��ұHL|�C��>�Z�O�*�lZ`�&Z+} ��M���b��]�иK5�+����QX��Ƣ6�]S���C�"��#90Ƭ��8�7����ۜ�}@�V5 ���+��@a�C0�F�Lǐ���b���E�je�d9�ᇛa�nyw�^mxW4s��
G�X��Rh��Gǉ������R������eC ����+4�}��gd�L��" ����e8�m��/�����A@q����`	M�Ў���҉*&�Rk�urq@T�t3,#_͵��辬27(!��F����kxE����q�L���g�;Y1C���DԘ�K��t �S��QϓD�)krl�Yo��m!0��V�@���`����l}݀�����O�����4a�~=�ݫ��b���/�jq��63�E����A�Ǚ�����%ŏ��3�L��1�C���6S��d����}yoOc��@�c���SH<f��A�����ץ�\B]J1P$D���&:b�:��Zf�h��k!0�(�G��/����h��3�Py��d��Ļr	�����;	VQe�
/#2�85��x�2�T�x��NE��#�:��I�����J��"�p��QH�-�dlO�V�a�U�C����8���e&��`j�O>��`���ڰ��݄�q+�A43/��zY4��翡� .*��Ö�A�B�2�ԇ�6��(m}]U�;�E�V@Z��.���{��Y��;�3�5����͓�մ�q3_M=-~����zJ�I�d���D��3D�I�B�I�?G6b	�`��#,-Dw��D$�����Wp��5nP���1����	�1��b�K��8�Qvx���r����"������G]�,��A�H,�N�d�,��D#��+��.��6�f���73آK�ó��W�����?�%��U��$��������^�X
�y���&2Ͳ��ߍ�R�(�i"����;fH��"�;q��cxQ�6�e����H�T���)1��:Q��B����L4�"�iz����¶� �<��.�"�7xݿ:�	�B5�-��#����#v���w��c\f�^�c��K�/�!�"��!Ҏ�o7���J����ȨK|{Rӿ��E� ����$;^���,?�mѮ��Gf��"Ȯm�"Ag����������:)��S%�PmR�%BD���E�>��Z�z�x�́J���h������nƮ�B)4]w�&�����:��"������w�%&~d9�n�b��IZ2�.��zT
l�az7��0Bϩ��sr�#i����Y;�!��M�h\����j�ʆ�=alVQ��Sӷ,��D����T-������:R��d�Ex~���U&�r����kip�afA�b)�8��]D��O������s�z91�Q���nX��\PA��&J��Aa���ͼa_S��^5�~��*qY�Ͳ
Q�.��]]İ�3��D���ʍ=e��<hR�\������6��a�O]7J6ު�l�U��JI I�I�����%�;v�����u!��5�g�L��m0R����$���H;b
T`��y��r�΂N�p�TVa����*�o^��98��bJL(}�E�0�l�k�^�鷙@�_�c�����q[4���J�C���	J�(��wd�Y����	��N=���.�8|���K/r��.S���	qr��s�ؒn��f�WC?���tWBtr�|���|��-��s�������@N�)y\śѶ>�VF�I�Ԍ���o�.-n��t�n)jb�ˉF]a�^���E�.�Kh�����TI-�y�	���F'�?R���_wv3�����|T.�!��T�>�YgBsaV�����pF��(=�U�+o�F�50���}�35��&���<N���� gDgʎeNx#�Js}�7�$Ę�Ht���R	��R{ʸ��W�BV'�3�[P���Qy���8x{՛��0��%2�0��^h�`[΄����+��|�JڻC���������H�;�.��5X%I!�?o*(�LF=��'�P����ȯ��߆ÄҖ��	�w�:MIE��P0�G�ڇ�uj(>,��B#��}l�q���'qS=!%y�c���ky:�~+�T��
L�Y��{ɻ�d�����0Z��	�aƨ�0��s\�H�\{��H
+�#~�j����щC�<Zu`�����2���������t$��&՘2(�ǙT7�YO=��A+fr�Z�A��^�,&J�@�(]�����F{�Q�_��^{��*����0��렴�UHR���}��%�!1�n�lO��`|�I�5�&wK��L<8�ay��"ٞ� ��E��(D��� C�{�Tzyc����4~�*��z�kbo�v$]�x��w~m��G*��.�x8m
�ǭb�nC_5����!�gy��9|:� ^gʹ��6ieo�4�M�&��)P�A����ֳ�j��5$#I����,�@W*���<3 1����	Q���wɢȾ�6�ّ{E�2��m
����/��+�xKǞ�=��ZI�����K.L�Mϩ����,�"��S�R&Va�Y˴��1��P���-_lV"cy5�GL��C�`B���5=���w��3����~N����Y��;������Y_� )�����$F��N�s�@$�#��&��W^S�s6�t��2���wv���!��Ga��7�u�F�pG�~YZn`�����E�)�)��4Ly�G1�3V�/����eU\�E��k	��?���e�W�
����W�5:R�.Au���D��?��~������1
?���liq(@d4��3�߄^ ����y�����TZP�����E5&fӹ����d��4]2�3��>L�v0i,��`CO�d	�����&�*��g(��Jn^6ó��c.*/���r.��l�;h��9,z�[�h�%`ݐ�\m^�/�3(�-��*Ψ�H-���T�G�a6�i+$��#�7��v.{� V���勇R��M��- ,{��6sKn���ґ��D��O�v��D.#܈&�k���0rL$��/m1����e���\�3��Ŀ)~	����۹[�ͱ;C�8�t�FuW1/�C{���&��x��
�k���Le��~_|���n����3�Ռ��t���9�/�f��K��"_����kL��"�5�`�i�F��&�;�p�W��k���b��h]�����٨�7۵;���3&��"M�JLV�i�_እ��V��M��{��Ew9es��Zz�[�߂²�F6 �����H۞�V�,�ezt,u@9�9�a�.�C�
e-]�}J'�	ֲ��>�l�l�q��s�$����RU����?��B��r7��,A��[P�	�5��� �78�ɔ��f�D�f����i�L�������-d��408+c�y�&�0���$6���=��i搄��i`�o�4P&�F3!}DP"S�峪\���}bOG�Ġ����kd��x|�ʶS���ᬮE�>}F�*����O�i[�M^���9'i08�Y����`�?27辿l= '*y�Kcu��⇧��S�F���W�ǻ��2��ס��Q	Ѧ⊪�X_���F���|��T�7j�Vc�恟M[q����c�$��԰L�ŭ�4�/����*�:���ɇl�\�+0��x��Ŋ�ðU?y1PS=�w��)(S|�Aѓ Pm�Q�0�C�Dq~�Y��	0e]"�l�6SL� ��ks/����(�
�xv�T����K/q 	�� לr��'t��x�HW
 N�TF���X!�_���	�����~`=���eqj�����k�����W��0���g8P�/K��f"[>]C�s�9]�%i*B�=` Ȁ��������,~�՝�	A�9���o�E;�ɰ -�3Ս��/�z`<��L����އT����q8\���vR�l^=��ʾ,���3��5��߾s�>���]h��hV�D�Fb����jwN�?�ɰ�(��-WWbN����Ex�����1̣hR�˃�vc�䝹/G:��x��Ȑ�LE��
�Σ
O�ٺ��+�ӰMȉʤPc�o�b
�뻝K:��_�,�=��[�w�Bãۈ��o����m{?Ե`�T�Gʡ���&R$E�:td�Ib5�L�|�������	щ&'tס+{l�U������-;a�ߴ�)7���7l,l"B����[��/E%���E��+Q-���?���lk$T3��������6��������c"!I�<S�A
˪WM���GBۡ�~5[���!L�>Kز��� s�����Gk�jS��u���øk㛮���T���G1q$ɱ��=LN0n�-��9~�?� �+�[����	=Me��8Vw����A:�$��=�3�<,Oם�j��K�z�ݩu+��)C�_%@/o�#*��_���,�<,���g(�St2��@�����o�L���5�-ר1�j�W��$��S�������L���x�s@�Cj;fCk=r�VP��X!�x�h�vUK�"�8���"����
7��T�Uq8X���\�NK�[�٠B���bJC����I�m��"��*�ℹ�8`t��"r꿎��l�z�(F##L����`�bm��>�����j�5y�P}���Kzǈs:���7�I���]�b&���`ү�M�A��ji<S��v�ꨂ��~Nق�ML��}�.u�i[��t���Uz
'��yZKM��Y�"���d���S.L%�Q���:7�NG�4��P(�x����������[�`�O<�f���N8a|���%iֻw����E�6��bg����f�<��N%l�W߇D,`��3s.ϥ�<��M82Y��+�:��'�ż����gNN��V�*�4"o&P6��}EZ��@Lpf�Q踇�� 2����[ �y�d�����
}��x��-�(!3:��:��+�ɿ��+��zX1���$<(�ۺ�����:��_��Y�`�h�)�u	���|�k���v��?A~����)l�YD&���O��BF�r�*"9�$+fR��,3�e���kS�#S���~I�UgAD]X?H�&�_�.&�cFÙԒɑ�����\J��nTW��r,gZcoY���R�3h�cF~+<B1`q�\W:,����U�`3�)��'�Z˕>b���f��e�h����O��/m��1��JpK{WJU�f����u:8*���u�?�^&���v�����3���d��xe����[�������ث��s"����jA�Y��\0�P��Dz(�B�-sݫ�!-�=����ݝ�Rw_��Ֆ�#K�`dZ�G&qF_���ATfkb~��o��v\^D���骵��qSI*O����h�*Eڝ/�~�W�'>�|��Hx�@��������n�t���/�D����u/헟�o��hk��dL7uη��D57X�?mI���,U��M��g��F��0QJ݆�Ύ�5����hs}������PƵF�	����$j�������eB�q��x�	�
K��8`YLcT��3!��u�ݙR��+K����+�)�����z�*��s��O)I�/5d�C�vr&�Fv��k����v�@3Ӂ(��`[��8B��`���m��kj�D�V��5z�N��m�"�h�9� ������>���@u�E�z1=��[�?!��[��B��6L�8�#AkE I^�|:���Z� X���0���j�.��1��碅�y7:�n|,���)�Ù�&z��?�I�����*o8����]����ˇ�;��ű#��*�5`Z�ZH��[��^9��'�)U�{cG�T�����e��7�Gf0XJ��=�,��x��_Ħ28�$�a���"����A1�Ye�r6����֢�k��@;��4���U�Δ#�9	:rm������������	�F�|���&{��rD\b�.T���:uc�U�\9�]y�[Pq;4��Gb#�W���Í�t�D~��of,'�!��J��yY�7��/�|U<���y�0FHt�1�˚ �ފ�xU�()1��/HB��ݳ�\����� ��	����9!���hbU:�h�1YD/:[�N���E��ӈ�:�J�Tdg����T*
��M���2�1�B����:�����s��nz����������jo<�r�.LL�"8�뼏����G�Mb�IR8H��m**�[��4�ݕւ�3Oi��r���"_jFl��f ����ϝ��-�|lZ?�C*y�� @G�ӽ�cH�,B�w�� k�S�.'7�h���`�z�%吓���2CD<\E�\�8�,����+i���yKܯ����чf��D�tu�o��S���|�T֖��ÄEe�R:*��nm�`��{DDZ��
�uz����򗨅�i#^��*����R�a��uv��'9�l5��;��kϮ�8��T�zM^�_Hu(�j<�Z�cJ�ml[�|G(��h�"{#TwqR3G��ztﵦ����`�G���WF_�/�w��e`O�Ķ�����$3��@���d_� �����pp�tW;��w���s����'��r���j�۫���q DA�<��}E�ς���iO�C7A�'�u"�G�_S٧S9�B����-�C�/��·uk�
��Cp�*S8�d���1m�u\��q�PL���~�hz)1��XF�حx3��n)��pRظ��8U�,?�����@������<"���gW��E,�X1\b�|jƇr>�G?�=o�r�k'vjؐW��6�=�w�ma
6@]��P{�K!��N�����C� �U�;�v�ܶ��� R��#�?�G]'�����b�0�����ʜ�B��]5o�v�M i�X�P�ȝ�.�
{��(���]�!I�&y'Z�ʞ��]��j#/tc����
Oh�Ed��"��o��\����6����g�Wȼ3����B�o�9�mc�c;0L���B��J^�S��t��r-���wb�������/C��)㮹�Ϊ�(L ���C��o��tl�^���yO�I������e�.#����S�+F�ZA^<���_x�P��R�'��U"�@ݔ�(�ޥ���@��Θa�`a[J^�ģ1\[��@�����-4�F�J����ѐ�����jH��N"n.#�]vv�2������v���l����2��[�ک�O����r�����lT-���BO��/��aX���;�DI���桛����S��圼K�ʶ{=eQ \
\��h��3���'z�vp�w�Mj��טQ��
�y�?%_��v��i�'���C�%a�u0�|=��Y�,�,J����#��}�9���kV��
����ƫ�,�S=�!XfS�$w0�+d��٣�oFWE�c�FÔ@A�L�Zl�*����j���b�˻^.�V�~]�yw�<�PWB�{di�*9�)4�ǀ�T����C�od1�۞-<�|�G�`�~�2�>�
��X�����̎?�:�E'1����P��4���Z]m!���A����U��1������}g��Eu�j���%'�Ɠv���]� �7���_�җص�^��\����I�LN�^䊤��{tn�Ɇ��#��6q��3L��:��8}ï�W�P"� �1Z�3P/UYO���i=�(�my�� r�>�J��m��E6|GI��2�G��3g&0�.��O���FnW�ڼJ�� J��M��c�3O\��;:3��qǣCq�t,梿�rbԘ ��Itx�悵��l�� "�pn���"�z �|���{�BJ� 2N��Ss�î}�P���7;F��MhB�P�JQ���� �J����Y���u�;��5�����n��f�>���n�-(�8�ð�m��yz��#�IkǊ�n5�m Ŝ&zL��7� lϿ���ʩ䬯��S�����u?b"_���<�X �X!{jA��,��� ϩ�\��z�M�PnJlL��4��J�&#|��N������aO���r�5�a��3����rC�		�]ʟ��q�A�,�}���^gz�s���@(J1NIV�q��W	ự��"�%����6&��XG�Y�L�����H��\oq+X�w�':��G�q�.��.=w��`昦�
�'�'�T.�B(fb�Z2���4�^Lu'���B)Ǚ, ڿ�Q�gz�(�8��-�sLڲ+��p7���ū$�O����
��!0��=��iv��x���+~�VR�k��s�wW���~M���'���[*��k"+h��G��Q�kg�W0����Z�VM����&Ջ��,O�
5^�\�r�
��ޛ��~]�=�L��I�',zi�5RtW��l`L�X ,S���>Lz��;�T?[:����M�n��Rw3&Ew���z�$����!�>�<&�+�^R
�'zyO�	/q��sn'cL��<���u��yd��! !a7hb����8��u� ���ա8"/&��4!b�8�fQ��,���XlFt���f6��4�)�8N�
n�C��ԥ�E��S�k�.�t�p���Q8Q�a�v��V�L�9�-s����Z�q#���I�b����"�KI龨8კ�k�2)W���r�#�Ps�(12���
��[�eS%bRƌ�������B����aQ�i���$N�C�	2B��=��S�d>�S�]�eq�S���߿|����Ι�rv�YVGG ҁ���z�O%v�ȑ���1+C%z�]$��K���F���k�RŌ	p4�|�o�J�4�d��0���i�	#�C���
�C��*�1�lw�.�l-D慹T]���*���˷�9�1��U�tz=NM����[�����$�E���ڙ ~�Þz���\f���R��K�e~C��@�2�����i���ä+A$�7Gr��l����t��DD
|;���W�-�q!"T-y�<� =D����觷cN�"�a7����\��&�҅B�0A�W﻾�/�R��e����Cُp��D�Ğ� ;��}T]�W�@�j������O� ��U������*@����u�&p�4q�+>J�*���P�l���D]�����&�γ�����瀾�ZP����h|��:�F�cWux�����1�ٶwi��V+Wqf�t4!|��*��r�K��� ��&ZQ��̦��	̈n}�_��i1�2��B�f7[�
ع���-A
��q��?j]1ݪ�=��!���Pvg$t��{M
�����05�H��I,��]��af�	�b�Q���P����}��>|\P
�V�Zҽ]x�I,B�DN�;ғ��5�8�����/i�T��>��70G�*a�:a
jѓs�������o0~��"��~�D�_���>-@����W��β'n�;B��5�<T��g��@zM���T �ʣn1$4��>M�/g�H�6�ك�^*>B�g��t��{ʺr_�=�bٰ>ǸZÈ3�3˱/o�-�\3���vd�R���d�4�]�+������3-0�9��P�1������fZx��>�k��'1���1����h�W�7���YD6\`|\���Zt4�mX�������>�S�F��i�+���E�����br�z�Z{�U��X���se��Z�q�m��c��*y�t�����-�CU�#f*��~l:���J�, qz�=	dE���}/�c〙�#���L�z�z�(J-�5�e�op%��s�6���D����cFdh��иv��6|��9-�/�R��ԫ�Ft�| �m�� o�b�j��˗U'x�GÑ{�G�O�}I�;o�'wq�A}7�P�:���e�����ī����,'h�v�_��?���̖n@��{lR��]d�jv��+֞��,�����fv�����w�����z&��k}���Q����X@�' �ez����^A�%���	�Hk�*��T��o[��"CͿ<�<��
�c1�/�'�p���>q<v�ضu�����V/�0�&���B]$������-1�؎���z���)���[<z'�{;qܿ�3d��0d�m:�;�� �h6�w¦�u!h��<)8Q��H�>7���d
��^��"��?{/g�00���D�]�Ln�q�P�ѷ���7���g�G:�Q1�#w����T6K'�d7N���3
Y��}tcTW�Mv'�cڼ�S6$���f��O�4�+����d��k����ZXǪ�g����;0~z-~D���v�?:�ј����a�Y��o�G���P��S՗݌zdp����f���!n��[��E$��OC��<q{�K�wq�_���T�%���@��ye��m��,p|�_R��p�d�Lu�Q>�ة�וu�ɾ;��\ߧ�R���Ҿ�~��	�;�I7 �<<Jc9!�w���O�l8�aLS˖!
b�@�#-V*e#�������f������� '"�i�W�5�ZøJI/��+�f�5�S�O��U�q�+�p����i��p�#Q}��u�r��%�z��7<�����Վ&�9�j����x�w�ȗ���NjP��z�?D��P!���@�����Y]ƤM��΍�#-�kd*�ڵ�Txl�e�UQ�B&�����7�*�O��T���t:E;+i~��e�g"^�������*���d=����8@o��E���x����=�$Ӿ��|k�3���ǅ�:�d)M��]�ʮ��B0�_SoO��~ϳ�R�ߔ{4�bD�!Nkv�c�U�$�f�����Q��AZLz��	� ����&����Z=�v��n0�"�t�n��ʴL-!�/)aIr��B�k^�; �x�G�<�,��:A�����A~!F+�bp�����2�.禰.hix�����a tKG����G�BTB&���[!GD�3��S͓�j���#Є:����
��
W��n˟<�s�c��d�<BtS��w����D=�F�U�k�dd�v�!AJ�ǅ�U��#��+G?,�k��Y�-�
eԓ���`��t4fQh�d;���8�����":e��5�Fi���7>���u���'g3e���a���h��B5Ƃ� � T��E4u��ᒴ2�UN�4��A�SP�V~�t0$Btk��B���g��߇v��Bk���͐�Oz�j�U�2��>�����������T���9_g���N��#��A+N𖐦�?�η6�s3d��]rךv�Y���,�aN�?�bs6��f��$�,2#{\����#��p6����d}Ux����C��	����ċ�����d�c���4�g��PzrY'���p�oH��X���n�wV�Z���l�^�B�|\F8C�E�P������i��.��sg����J9'?�/����·k�-���!�0O��Y7�5@� i]}&P��uYԷ�k�}�h�y|EM�)�Sc��:�%o��w�K]����&p.�r�5W+������C�'e�w�A+5�+�fȋp��hu^��Gq�Cˁꝃ��{a�Uyw.���x�LR�{K8(u϶B�T>�����1�T��nݚ{���U��歞�!�N.T��\�� 4�Ѫ\�u��(��i�[�r����� ������|g3I��%D�ZJ���
�mr�4F]��jh���S4�D<h��Ys���k���k�縩}fͦ�@h�?�5Ľ|lC���_�6���qR�SV�c�.܈����dd��2�����N���T>����'�/���~��֜�K�����Þe�ߚ���]�[
b��<�qS�[�D�.����c�`W��@=��/�^�P�Q���!2�G}�	x�#��8ۺZ��æ��f!)�,�<�7&����;�|����**:n- E�`��Nk�lTrˡ�_u"�#��PV,i�`u��WWA�I��A{��3XH�8S�l&�f=u�V�[=l4�7�@`T�
�i*���EK,�`��˯�f�z])m-��r[ຈ��,Ii��C2ؕ�v#��V��S���#�SZ)�L�a�1F�u���x�^y�&3a��_��zf��̿L/ly`V���3���a���R����~r9�Pư�1�ȑ:5�$>M�����������%C�Rt�����T�S@e�ғU��7mW+��J�z��s��i,s�����I���|�Dx]y"�]#	pU^|�2�ƒR.��['�k�����6)�P�ꛔEAo����T����/�Z��M��ٖJ����
�+Rw)C��#�ϊ����YO�o��"k9xEU��u�w��?.3�>��#�5���9�)2�[�U׮ļ]���k�7����;�Ŋ���&6�}���m lo˨�&��.���У{L�.��n�Ny����1�tطD��{~7�%�{Ĳ��0��v��`n�iU�~LP`fFa�G,�������N�!g�Ө�{�� ݱ���}��)qc)p����
���q�$��^;J�-�arQ��6���cՑs]yn�=�Rh[�)�}?�O�0wn�1�=�Z�H0�3�?������M�:R�7���������1+�XQF

�S�=��\�sPN�41���)���ǌ��f9������oA�M��8�椖w%�{�M���,\b��k�#�э��n���'#V����#�`PC� ;E�7�8!�]���4�D����ѣż�Χq��I��!��,���V3�*�>[!F�y������OG�ub}�* o��˱�i)�:�����{)S��`mP�7����/lʰ�»z,�������`ꇿ��Uz'4���@���^����9yyɿ�<V�-(�PSD%��Ԧ�r�&���������b<��b�s�O_`/E�G���e~�(,u8���3(��s���ެS�MN��#�>_�x �ղ��w �<Z��u����*W��"�2�������/=�5�mx�JP���X�C��+8�_�%�Q�VQV����kke�w:!	���
�eό5j����Gw)���+�1��;���
-$�xk�0�U�X�J�UU/�zU��C4��rT!\܅7��:�VV�m�
� �AX5�����_%e�y��^����wy&~��;'<��{)�:�quT.��=8�ˋ�W@��j���1��~��xf��2S3C�т��!�PWF��:�^q�^�N�I����^P��ܠ쟋��]��=t����:�B2��!��A��˖?�e�W�<.�A��/�Q�Oј���7p
�����n@�<�k,p��g����RZ�Ү��e��v��U�� �zA��%_�䆏8P
ᬫ>2���K���J�p#WsX!V�t�q�+�f9���t����Z�>M���~�պ�E��2��o(9$�6�BX�q��n3�#G��g�����NP�&d���%�|b��?~F�"�h�5��#/��J' ���4�+l��e�� ��Q�0]ᛀ�$ڜT���L#���S �M��
mfz�C��05+��?���k��-��n\���ڪ��b����������)˶v�_D��q9�1����p�4��P��ˢ`I~l?��Ƭ���>�|j~eh�F�-Q��RJ�jza�>�1������~���6���K�Kl������2�q[,_mN� V�]"�N[�ͬ���?U���;�z~#�}��p�%B���I�Nj�4��cǆ�l�ahNu~�����9vx{)=t�,x� !���Гzqfe�>yZj t�C3��~[g�u�v�$�܇;�3)������b�`����hGI��n��RB�M�`#Z��޿��(jv��%j����ˎ$4)�od�eh]�i�Q�M1ƥRdP+j�
���:GZ0s������I��{\��k���Qp��7���I�FMo���=W�Ǽ�=���M�{O�L0�$$�+i46����?�rm߿uJ@���r�^�D!v���6	�,V��|n�^��~�-(�T���%�;1�W��Qꭒ�wy(�GR�h�,�uƨ���|?���ȸ�j��+Ŷ����x��aT|�,��>a��t2�ю��H�N�S[^�)�4P��?m���|DXI]A���K-��_am0�c��<U��;Y�nސue��I��'����D�;�D�rF�P��`�/�a��a�3㍠v%%E�NpF��k���~J������(���%\���dKrj��d���\�j�a� ؜z�&���實Q��P[:�� U�{���@7�[�wX�˱�L!�ԉ�x�97c����P��[$���tP���m����܌d_#�5ύ��7/Y�nu'R6�V��2I ku�A�I~���+�+���4�=�14�4V$($��v��E|��&�!�x��$c@�gGw�2	�q�
3�a��M���R'�c�k׶�F���*o���l�����xqK���[r!�:l�Nę6F�4R�"X�@J�J_J��4���{�=hӦ� ֒b���3,#Q�� ������w|�	$�WC�'�`+����Bʖ�#�-�`��M�F|�BO�^v�?���w+)| hz2�9��}�F�INUw����uB;��Rh!�k�6q���H|�Wŧ#I�L4-2����}W?N�-tƍ��Ճy�g��%���)p���y��ސ�����ې�E���"�p|��f�Hb%bTZ�Gdq��.�f�ҽ�ֳ.�+<B:d���E����Ⱥu?����?"˨= 1X�yy�~>=��R��NQ�P�E�� �������������6�i��
��B߫����hȺ�T�Ўi�Vj���Sikv����P6���G�}��"�_/+��{�a�[�r�A�\|=��9���X~V�����>U�Q���R|sc�q�D1��?�4��04�i/��Q$������zƀFw�Kd)2��}��?�n��CL$��
�D�]�����r�s�z4hp�g���3RëR���ٳ1�o���W8�E�6�T����ި�e��ZԽ��J&Wbi���w�+����؝�'Y^�PtA��C��ωGC�����`Y��NʨHh�9F��/mc�H=�J��w"��!2�I@L�7C>P�ڗ�C�uo���V�b;3f_���'�i��MEvff~��� -��6�����jA�S���ɣ�ڔ�k��I��v�ܬa�Α|Ы����h�9t���ZͶt�#�9�@���L���./�ܓD�0��ڒ�$�"�G��^
U��R�3e5�h���)�6���"p+;�[��jB��t��xӸ�kF���Ya�a����H���d��҃SǺ<���^qJs�x���5�U�'6Y�����@�3"-��hۗO⩊XI?зo*������Z�EP$$Zkܱ����^���Qi�v޼�?�`��9�i�GO�q�="L㈮�ƚ��Hz�3GFL�+A������2�\���Z��Ƀ���޼o���4��rt`fo�ubA����<v�pծ��}�p?��yŕ��W.�A�ǭ� teW'_��gWD�&1#�9���`��� E<ELW�^���w��^͊I!L'���?��@���S��O�P?nV�c\�Q�!g��ơU��Q��Lv^twCW������P0!=[�̸=4`/�P��>Ҝ�&��	A��ot��PS�u��됂TE�v�p�dA���iτ9�������D8�Q�X�u/R�H�4�{��]��ܟBlJ�6���w�91v��6����`�4' �W��Z7rԃq� 5���謰O�9�g1��)�7����3	DatDDS�{h�׮�������e�$�2'���cX\0���M�X1��%}�B���/=���x�EaN�˂�rp4��}��t3V�o�;w6���"�+S&����)+��g^�W1Z�4�?���E+bD����CG���і���W�
[�A& ���?�Y0�ï����=ϯ��!烂A^��/2�H�rh�m�i1u~a������j��S=5b ��@~�^��e��2~+Pܑ�C^�(��}�a��Gi-.����E�ۨam5��m�k�p-z�b�n�H�-0�~���跏����ue�<#9¦�R�eh	��Q�3Y82#�Nݜ���oUt�T]4n�
~�6�J�`�_FI�˱�1�&� �Ow�Cmt~6���r����!vf�V:N��DX������T��J�̄d��A*x�C�� ?�t��2Vl�buD����G��z�byH�V2�;��W��fQ�U�ˌ�e� l�}�J�p �����wC��bXxů�=��G+}�#�3�s�5�|�|.t�O&V�\Z̵Y%��$�'p\l��n֝�b���wC�S���WY�.�Х�8��X�7��v)��C�^k�U�xA&K~���$[�a�n-�P�Q���x'�1���� %|��k��������n.���k��N��	~�i�?<����,.+��6�kN�g��� F2�*����nޠ��<Y���pB͙4.T�^N���	�����_#�)�Fd���&��Vvc v����Ll��)e�<��|��:����T�GH7|���OgyɐW�*�X$�&�T�P<�"��j�����?�U�CݗK���x�n��3��8M���Dv0u>E:�&;.�7�+n�Y�z�) �S<^6�PC��#uRb�b�"�h�m �	C�z8���BϖNvu�1�mZF#�ث���D�y-��~YΠ�����N,M���f3/r������cA��ǈoj5���
�����0��cƕ�pz�khd)�,�&�=���*t�RqАz�&�<��3����٘у"��͛����&H��L���2��N9"QS��i���ydd�y� q%�	0!Q7��٬)q���G�d8WI���No�`����6�S��|�/��{�T�zL�ˈ�Ce?Q��yչ�X#�5vM�
���s� �O�y�ヺI���lB�m�j��z�\����m�,����������� ���:]��S��2���?È��XW!�/娊��,0�^�LE�!ʄr�d����K!�]'܁y��{�8
�o���#�w����ہxǱ�|�֒i��U5�@��٥uk�Y^R_�FM��]�7S�؅#Uyxd����O90��0'��U��J�2��/��"���N��������AX8�����j��SU1����y:��I���
����) �q�}��0���$1Oa����$g����NY����(��Ў�eBa��ۃ�~�J�4#��������%ă����Q7j�(n��yp�9 �4'�p��͎Q�֮g��<ϐEG�{<�b�5wP��Gy&v#�hX);�Ǐ���9�f��_"�[v��I��MؼIĮ���`���*"�lp�5�F=�����!��qgխ4�7��
�{G%ց�)�Ne8�w�/8����@6[f����9� ��L�_�ͺt�H<^¨��W��zV1%���R}�aӤ?o�숯��Z��@��e]�Rs��KO�s����T]��A31[�MU��D2��H]�5���~@��׼�e��[X���^ٯ�������B�J�W�pm&|p��q�:�#v��TP�HZH��a��+G��l��`�C1)`<ڇY�K=q����4��_�����#�R�d2̛}�F�nS�0
�3Mθ��f��*Ԩ���;�6�:���y����rT�3
 A�[n�b�42�?�e�t]���L�.��6q�}���1\�]��7�� t���uC�����R~���p�D��e-���G�-�3J�y�׸iAW���Szq�j3ȵ٪|2�L��:�&C��q�����mfPڻ=�8s�����T��C�[
+��'�8��CV���6�� UШ�lz]�8�2�" k���Dg����T�T���>�hY9&͟җ3d>R����qi���b?W�C_/�FU@��p��[�@s1�ة')�A�>�����̂�yn�V}�����j�S4��eD"����2D��wq�D����؇l^������)��8y3�Z���E����/SG՞�"
�*( ã[��&��=4x�4yċZ[��bO�ٲI�]wP롴J�|R�yFoE��U3ȓ�M�j��E�.��JU^pN(�"��_�x'��P%(�J�����+A�k{�w`�9&˅����˵�����9���ľ�碸ʢ3����ko��B� u���9���5~b���`uY]B�l���x3@xI;�E/�����q��F���ۏ7��ٟ��iOj�sS!`C�i��*	P�2nH~��������t���#by��qc����|=G~Y��X�Z����q�C��`G�}����Oƕ론6��ˆ�o�>�����^���f�Qx�>�)�>e��R�ph����� e��4V��cX������uZ��ٺ���"-��Cߍ�rv��ڃo��՘|I+G����x��=�X�T�d��ȶ>fK\�����q�ș�ׇ�4�+{���mV������������~ӂ%�Z)���ؚ��aD���{2�,�u,r�G��?I{�O���~h�����@c��l�5<U���A_0ƌy�C�lK�,�r��l�J:°ә"F���`���6�9�W�~?l����v��อ��Ne�xR�zǶ閜��+[:�z<�� �_
O�H������j�3w�C��&ް�@���O��R���/NOg8��*dO�8r�׳�`��)��R��!�����	�{�p��ɷ��˯Lq-�c�Y�S��V͡��X.��J�D�k�ѯj~u�t����{+���� h�T���@�~k�ئ���+�������ɧ�wr���P8L�v�bF 	,xm��Ds-�qM<Ҙ�.���SE�L��n��q����>���K8t���{��Dx�pf���'��i��#rlp�
��b�� ��P�a��{لKOZ�#j2k�{狫h���|��R���i �������w��ItL�M`Ks*s<�b�Ҷ:�<1X��1H� z�k�LTr�d�~��}0@�v��}놪������K�~5+��>;R�֙�*�c�i���*nQ���[q_�";��T©�Jy�R�L
�Pm���TF<�7���~Qy	�����Vb'����^�qe�EDƷ̉���i���9��u�Y����)[L�ծP{��˟�8��1��XtTKjä�s7q���nz7�_�y*d*�M@���5���@� k��;�/��޶<ײRE��`רD�uH0ʌ$�u�?Ч�gv�d ^�~nzq���L����谄�YE��oׁx�a�P����8���s�q-�1ϛ�q��m ͘�c7��S���w�������Ѝ��ڻ����$��x�>��H���8���Jb�m���},�'@�%[�r����5K�]��+�Ʉ�"o>��A����O��\z|���F�̱�> ��~� Ve���Sj|h�X�����T��q_ ޒ��~���j��BϷ:BW_"�k�Sua�(��b���5�D�������Tú�蝐��A	�A����^:��T�'TQ�<����n��crl��W�pQ�i}��:ͣ�Z�W��K8W�şV0*ח�?L=m�s ��ۢ�I��ehG~�����Q�4���an���@�]Z����b�E�m��RU
w������@�8�}ۨ���[�ឬ��8p���-=c�M��h�L-ﻚ	]���������D+ǖ.�*�_�@/���{�Y`�������w�<x �C��P���]ml�ol�a2�ґ"٣�s�Wj�ŀ�&���W
��q��,)4?ôL����w��i]s+���AE� C׽�	:^��b��tm_w�����U��R���:X���3!D�3�a{!7"-~DΚ��;|�	7��G��t����}$��~E�E��G�at~N{�n�h�#Q
�����:�l�����;
]$`D_h���,3J�Y��K�����$����/����m�h�`�1WlO������TR���U"<xyzMQf��3Ɔ}P`(�,<7`�n�0�Ϙ�"�g�M�-�uC�,���i8W~��+��%�ui�_�}��{��U>iϽ�tpT0������W�e�|�E���53
Z0�f�b.�����(�U��{�m Ok����&_����Ρ�׮�iV���V��Q���kj��T��ٺ�Ir=9�s���y��mZ�4βۀ���Q2ͪ|~��\�|���+UN�m�k���c�u'Y�,�1o�e|�sC�p����2N�I��8����i:P[�HȤP��6���Ij�I;�h��K4W�����~%Pi1�,��͵,c�*/kR׷��[��6��f�`4p��	5'��,B�[��ڇ�lBz^����2�i�l5:"�	��U�����D�{|���$!9oVD�HA������H���9��Y��]e��B/����s�B�[یs�B�r�--A@���_*��P_���ޭ��X�4���ڤ�;�\l�=�Fm�p�������g�0���!�z�X��ɸ� �V�Sq+)��{; �Hr5 ����n���xWިv[������W8��fn"4��I�Ű�|~�����}�TL��Us��+v��P�7�C����4�{.�7�4:X�+��d� ?��O���ۓ!M�Ӹ��V]S�)!�V�^~�ܞ���=@�Py� �b�ra^�M�S,6	#�0q���3�Z�m��S�cM�_i��D6��^Z�l�����&�#7����� i�Q �9?�O�6ݓ�t��g�s����
R���.� �a�,�)�D?u��B����w����E�*]M��Ɏ2&�]�+?	�����K��_Z6X�j2m��f�^�!��b��K.���I:���:�t��g��ᰱ�}���tpʫA�F�?��=%�x�K�U~g��LRR���a��?�r��*r�h@�/�+�(꽑54d~*���\窜|o7���24��B:������Cm<��L�y)�V4 >�ܫ�>Y�z��B���m����6�\�������3�u�ą %n������Z?%�;0'���=e�z˼&V�|�T�&��6���Ѷ��M���	�Ñ�rZ�!����Gw��t�$��'�֮�lj�;�_�K�i/檣G��a�.j�[)��dՆ����Z�� C���O���).�*��ʌ@�t�},��	@Wv�=dG7�]�\|2Pn����CԷ�=�8$����i..W*^���)�#$��0%��h�i�RINf���i�v��q�#Jm`�GUBZQa�j�n6b���Mv`En�E��\.�t|���ڟ�M͠�	� ���fI��H��ޢ�и���y�3�<��y��I�JP�i��J�V��,Ql�~�w���iŶ���8]�~ė�Ȇ6�HڪL�I���u�i݅���\���X$H��Qv�nٛ����X�0�-��_���F`7f�����\l� ">�{��iw�KQ�Ck�U�t�L�=l@�k .z�9��u~	#����ޯh|W�I.ͦ0^���E�
8(ML\�U��2e�A��ŭ�)��P)��	x����*�+t��LT��.�Ϭ���q2��hs\�&�֓�.gM�3��.,��78�� ��������(s�'Q��gS(L]*Yb��/���[�P3MBp�������s�0��OD�셖]9�k��A��Ĉ�;�O]� t_jϭ�&:�7Qd'QW�V哲8�L_}S�!N�J��ܺOc�	�����E��I\�9G��ڱ-�gn8��׏�a�d
4/e����;�ܲ��$m��Q��6��$���?H�0A����;��;�xo�=4^��hD5��Ȗ�����^gx7���8��	�:�eﶡ޶b�W��ͤ>S�&K��%����7-��4K���`��I��)����}�4�����:Ys�R��9�7��$�d��L�+��
�j�c�!��Ѵ��ZX��8cU��,E!��B���`�r��UKzJ�쫩-� �{C��=zm"��(
�Kr�]+%D��v�Jm�F�p*l	 lz+?�]eY�>�Tz�#8����$fis8��t��<���l�p����`Կq	��y ��-� ����. �+�g��PI����X�(�����bL���ʿc2K����oލ6�Sj�l.bXO�M�=sde�]<�@
���{�Q�FK��w A�'3�=7T�j8H"��7#���� ������*�'70�x
�Q���S����koK5��_X���M罥'0��$S�0��C2�6xW�[a'>�4��R���Nbo �?���h{@�xHy��q)�&X\�b��4R[�ßA��o׺2so���:�k(Dl�!��N���r��{=0aΕ�ٓ�������;.;�SL�Ӗ��Z��2&E)h!>��D��E=LI�&oH��.�B+y\_�|İ�^�!_JQo|jVz�M;�]��̾�X��Tԣ)\��U�������W��:X�����&�z�Q��G3wA����d��������PÞ�3<�
��2���	�9+
�]�'��w�.�Cؒ��[л�@lm|s�S��4��&mhF�s�����{��5�� �;�X��NLاFG_z�^���r�aӝ�URK>=�vq	W+\��:�ºwc�z]GWf�=
EX��	���Ш,�P�y�C�pe�<C��{N�E���&��]�O��`	�D�j��6��sjWC$ZĪ3��ɕ����r��5�����w@��Y�i�C��1�eԑ�tc�'�O�}�SM̸��+o��=�}@�x#Vt6�`=����e�~�6��ƒ�;�4b����|߮-��o�a�1JH����X�4
r-�~KK��X�T��	��$�|���,���~��0_��J���d��D��Ҩ�ǜԂ����q	��V����#P�H'j'@h�L5\��D/���CbZ���a�o*��}랄���JN��� ��f�IU�c�sk�U����T$𐓠��x�~�
,���?���'��)��	�Y3��8��*�F�gu���yw���F3��F���~���oJ�o�6UO�8��;qOBh�J�	��?��OC�l��F�a,S�s/Խ�� V�X
��2{����JhE���%�C��V5 �B",��x-ɢ�ZЋ�C�CO`�[x\n�X�y�At�1_�v
���Lg�'�'����O�t=_��6~�Ն�ud��3�t�	��R <�N&TQ醂�k����_ћ�Z����T�c�b8*x�&�I�BN��(s��Ď������?��ں�H_03���%��'�ڈ=���&!uo�Ҭx�+��;�8��T�휸��Q���4D��l__@�#��E�`�F1x�:7	�仅h"�M���,'|�MvM	G�S�h0%��'�d/�o%7���X��}X�6�=��3-:�P!b #�ĖMt�$x���o�wI�(��9�F�J��<F{�S�����:��?̇܊�����a��
��G��W-�ޫ��a=��a�z�3�ͬ�'�p>�l@��U��8����ވ��WB�֝��GНSi��h<�,�w}~��h��U0�})���Z�ósg=�C��$�l#.zP��G\ezS��$Qz�?��(��̿F��5}{ZO�z��8����Gf�!f�1��j,��h)���3%�W��0@<�飯���F/�;�6��ADYN��[���A�ɗ]D�
���NQgc�kŃUG��4�%k{)�ϯU0�i��!�?��r�b@��;m�|����h�ͫ��Q�DX#?��F;L_	�/��n�pm{�A�y����*�H�A֐�x$rG���x��KJ��,/�J-1j��G	���Ԕ�S�0� �1i6�"��%f�(�9_ m�p`#�E/=�r��ۺr��-�1۩z�Wr+��%������2�B�&ǁǑ��&�(uK
K�Q�E�wP��5�բ��S�cUڪ��<�� ΅8,�+'���z0�v_�� �����ƻx�|��?�ލ��d� ꝡ����#�I˱��3U�vh�Ƞ��pbS'�PlE�����H6;�lP<k=
�|D��)L#��j���,��+��Y��b!��(7���T��F�o
}N�#U�"��Y�v����IV[��1��{��x�и@�/h�!g2��6���/KB��W(.����(JRUC~J&���!6_
#�m���<nĄ��Z%䨉����?øHB㱥��¶�G��3BC�pPi>�8n�&�Ja�#kZ�tT���Oi�v�~V�m�"�\\9�H����Ȅ�����H�KE����`�v�����#|Z�3U�ͨI@M!2�|C1��"��)k ܒ�N��Fe�jgd���ǡo��*�A���ۺ|]�2���Y�����3�7W��⡾�DU�tcy��(��t����p���V�4������3�۴�R�)ƅ˭���E������� 
+�Q�XQ�z�T�L����H˩=}#�=���'���;?-�!���B'����v����E�#��8Z���z��v����#Lg)N�nJk/�7�a�����6_`@�>u�Cj7rc�FGS��^?��@+�k��XFx=ĉFحi��z$�0 ^��c���$�@���F9�w�,
��^�]��_�@���"�_S��e&���f��A�%: c��Z�2�̈́�_�}g�M/q\�t�D:������D9:Z�\X��eFA�![J��(��q��;g�톴����cb�%�{��Q �+^�����V�xO�ɣ�*�3�h�a�dL/�=������[x�Z�!��S���gt���)�~��Eoq���;�F:�Tֱ6$e��7�S����!�Vh�%�PE�	����'H.���]�v�����I�S��O�]]?������iJ_GsN� ��)a�Qr���'
���3!1T5+hLX,�r*��=q����F������oo����{j��K�5G��2�uO_�Q���"��h��T��wi�V	h��hoy��{�HT�p�n����QJ���a�f���O���ȉ2������!>o|�T��|��$�5^Zv����F��f�R��b%�h:���!E��a���78F�/Z���d!7��cC�.EO�lj1�K	5����7�k١���Qi
�,��J������/� f8��gT$��a�{�[��An���a8�DRuIJW��?`���Ԃc:[3e�'M� F*�$/K�p_���K�^_E�U����XY��lH�7,,m��	:�F`)�ɾ�k�� �a���:�u�:���J��p�\����H���!{�c(3!��?x'/G>w���|�TY��k������u���@�^�'٦�/z�R!�9�<j=,8�T�a�p�;7-�`K�@�w*�#�H�"�靠 4�\�4$�֕VYi��ݞ�c�ȏ&��Ԏ���ꈔ��U�{5��* n@
���u�O�~��c��ߒ�cY=o\.|��g!0%�a8����#�m汽����y��2B�Y
פ�E��U�h�h%��k���:V5)��)f2�`��>��11�v;�s?G�o��GyM� O��ȉbڀ�טǷ����*Q��3X�;U�}�:�A�֩es@ܤܷ����܄�N��XK��X�`���Yj��p
���;��(ߛ�>����d�2:>B���)�t:�����؀�RRD�1(�u�e�J�hv�/M�_m�ņ]���a�-�gj��Hwq��-���ݩ��3Gjr��"5*��Q�Ef�py���:�M�jmx\���������&�U槀����|���SX���7=t��m
� �������iA�T��Y)��oy+d��:��᮶�f}��=K|��!�=R2��6 �q5\hPL�f���@�5q�q��|~,_#�?u��)��g�\V5�UI*�y:S��^�xUޏB];%��7mg9�+�Wo�õg��ΫJ@�l�qoX�}Z��*�U�5̬�/X�ٹ.t�`0�v��Oq	BJY�A8BO� e9�|H+ﳰЙ�ʔk���_�tw�7W���L�.0r�~��P��˩��4��:Kξ7�{nvP��F����F��|��<0��N��/���0�\�\���?�����B�`C4)"�F E�{XCs�[��
��4ڮ6wP^|�(���I��t1һ�����S��hZ//�:b����87����p���_��L��I�S�j��g#"�I��!�I���[v^?"�M�Yߞ���b��_��=�S3�N�+��0�pA���v�;���?�j�=M,,��!���>c=V��i�1[�2��3,�~!�./�y�ѭ��W[S���;�~u�unh�)|�k&��P��b��'E��Jt�ѷw��F�UDs>j����i$���F_Jd�gby�gJ�*�&�Gʚ
��)��A:��e�Ofi�:��r����zڅ_��� ہ���V���{F��~�E����҆�H�U�Gx)"�P�pbwOB�;S�Gަ���i��R(�ÞVQ�W��
B���.>J�9����f����;�fdj�=�������0����7���lLe�J�Gj����-�Vh�i��!+Ƴ��r���
3�y���Ƞ)��bҙtS�H�:��dGO=ZX�}�������g��Ŷ�P��L���8�وK�wF$'��@s��<-�����ʍ{�_��řE�t��")'�N-^_e������ɫ�4����<z��
�	�����{J�9s+�v�]����03Z`f6�B�/��,�.��;��"ͣv��`e'aJΐ1n(�/�~f����&��o���NC�����rR�Zۭ���rk�^IPp�h!����1�U���S\�3�Xg�9t��dY�.J�#��i6���J�4OzH.T��|��ϲ�c��|��	K7)\Z����'m8|I�ln
�W�s�������q���������6�]�'�����Ep3��Ž��8��_��-���hB�����*�[7&�H;�;�O$$�ݒ˺ߤ~�UzYɂʣt>pwA`����kf�����H�1��Ȅ�"�s���vg�@�x��[��ﲤe2cf
5������P�S��G�_����`	ϔ#Q��P��v7�~}�j��Z'��.�9�
�}<>{�s�t�|�DV���N?��H�0�p���K7���]iBt'�:��	o�8��cbc�A�W6HG"yD��Կ1Xu<���"��e̕B��/G�.�$�+������[�B ��楊r�l��N��Su&u��a��W�f����)�[�DI��^o7K�9��m�K���];tV��ق ~�5�#�BY*��p�{�9�Bb�?ȅ�F��xoR�ɼ��{�N5���W��_no۳����HI�O�Jua����-��y��;�L���XA&�W�/���xG�u��=g���eݵ�9wak�v��֣�㻕�c�m	�Jūd�Ǘ]��V��Q�e��b�=><���&����>�`�D^s��tw�7U��_��@��x=�p�COi��S"Qf���ȃIy"��q�M�,��I(�|�7�b�F�$L�>� q6�+�'$)q�"S������<�ٜӳ�u��fc�W�aK��թWu�j����r#����ٰ���n�v�8
�Ic�]�P�����Q���E��2����"�7,��|Ξ�e4(xI��Eq�;{���r��zyi,���b�ɥ�9�\#<HD���C�Щ6��g�������a���sE+:l���Oy���x5��� ���~U�z����ə(�p 6f�t�1ѧ�DV���I��E+�GHR�偤<p�)Q���$�4�9�y����{���� �� G
]0����WX�^Ϫ��c�@~nu��/)�<dW~xyX��+w�2�=o'C?>�����MT�0����H��Zv�lrKO.��}3�P1,�0*Â�#�~�=��C�A����F�R�Og�9��p=ɮMiO ��yد f�j�=���Cۖd��T�\�)��_��f�K(`V5G[OVL	��?���3vH:�Ơ��.Fm�PT���
�ܰL�}��'���&C;f6��U���qBf�ںҙi�Y4tT���D_
�m�
2z�%"�(�e/���ֱ��oh��H��d��y	�l����]���-Q��Vů�6�Xi��С�.�2e?`P�a	l���`X���p4eamқ��su%�!{)���f���{0���ٕ!���_tA�mRH奴$�D�9��p�k2�ϝ+bN�<"�v�	�vա�YN���s��!)��:-o�*���9,6��j�B%@==ho��F&oGF�6�"�RS�kqyd��=	��0��`�~��VBw�=�`d�{z��4t��� n��ΜN��k�d�q�$Q]�1�^�g�֓DP*��s��];�͡<� �����W���_'�lm9e�wT�T�pfT/5m�޺�+�Ħ"����Z��✵5w
=������h-��/ܮ�=�n�*5b�5���>�u��LW'KV���I@7r��=2�d&��˹��`㈒=�o���ţ���x�K���2W^/��� �`��gq�L���t���>nX�Ȁ��|x�����w9��+���EO���ޮ��hdf�=x�#�u���he��s�B��|�c}�zdm�'d�+	�Y�q���.x��E�%]��/�?<A� ��W��t�1SZ��=;aܟ.�	��.��Y4r��>��Û(@�Nxͳ]G�`0�C����HU�:�M\�z��l	sU���%W?��G	ء�g�u�ǚ�}��<�_����~��	���&J����uv��<=���ʍ٬+)�d��$#�PCY�q@Fsu��$3	����%{����T���Ot�J�9|����a
�����iƸȒ{�tC
3�XZ�YDb�u�������D6�8)=txm:�Y�!3�TF�$P��3�����(�>eYQ��k)�����{ܸ�z�
�X��`UJ�Z�勡@��E�w[6��܆G@�J��H�$w>߶�gYx����:=��|0�w�q:�p,˭F��=��E��	Ϲ�9xG�MIPp��%����n~�p&G��o��)�)�|�j�"�V�r�7��U�o}��7�V#4���S.y�("7n���8��&����J��@�@�,޷�s�2�������,C�(K�,J��W�E�I@�k<[lK0��Zs%[C.e���~n�U6���qf�n��<q��G=\X'㿩]t����$DFjFc(`sG�PcA�U�$�y�}0.ُ�)SN(8?wԭt 3�G00���M�tV��n���6t̟*	a�Q1�%^��/G�'�g�P�:�mܔM�&*<�� u�k�S8�n�����(�s�y
��j����fo�.���ܳ��Wx�n���e���8纥XSWK��v�H�ᮾI�w���3��*!�cͷ�S���9M�\����":����ah^�R�^����-���u����\���Y��3TW]zBm�X�a�4%q
r	���*�t!�M/��4o/��Q#��zU�� C�)5E�cRw�E,2q�1R6���;X8oY�����yժ���m4��<��Z������(n�[,��S\�f����Ρ@"����3�y����n��+��-�(kh���R��#�z��Wg\(�"@s�k�m�*;�.鏱wpRZ��A��ժ�y� �
W�:�6�r�jP���v����7.��J��<bē�Q�soĎ�_�J~�6��vU���k��+B�,)k��#kȆ���(\)Ό�"Z��w��3t)��,��C���u�R���_��9��pw}����*-��E[V@<znҳ`��4�Z��坺o)��~c�;$&������c�n��a^���G�Ӯ ��Z0��WǸ��<�43!͟P�����ĕ��JbH�^�:ҹ�$ZU,z�.����W�e��"|U~@����,�@F�Wvx�d�"?�*�>Z��\��S��
�fU��ĭS�S:���c�²)I_ЕEI�7봚;����Ua;;��{l���[���՞_�(�#����+i&�ʥfk����nz�#:�3����x�
�T�7sj|�``0��I*)G��M�x-CJ#�D\nx4��L�^6����G�:� ��(cn�zMv����L�8;
������0|a�0����d�����t���� hK�&-
��2���f���	���7�\����q��@��!�
�G:����zON�/^��!+f#�����?�>[�PJh��Y��G��>�.�����x�F��/ )�lR>����&�w5((P%�'��n�Ō-���ъ:�	��G���=�a�	O�7'VlRk=f	3#;��[׉�5����I��Ү��z���bO4l�蚛^�[���\�h\�\&���4�`�׳��~p��	B�|��_m'a��8�m��8�)�P�Z��s�ߡ�ؓ��u)!ĊN譙pI��7]�l���4 ����g���r�D��eDH��b�2%�e�_U��C�mRy�k�ޫ��_�v݌)�V��4Xs���|;ׯǘ.|��p���A�*���$��q��w�?�2eH��y�Ә� �6N���Z�����������8y]�7,Y�����l�֑�&k�	w�.�%��}vdg�Ĳ�}FC�I��$�@7R���.ۚ&�DI�ʪ���J��G��;�ẃ����j�G�N�G�+պe�`��K��($�n�0]k-��ӓ��PI0���ӷ8���܍m����l������Ƕ��s6�\t�����Ut��\�e#qɝ'�$�c����x"��^�T��BTg9�6g�� ��DHI��������+\���R���N�$ߡR���\���/iBh���#&C����Z}-��lA@&�&8�uv?�w󶺑�y�R�)�Vܖ��7�d]v������D#~�yӮǃ[�j����`��Wyn�X�ݜd��M�9.y�r�G��a0�z�˹1g�F*�����K��E�s��7%�*J�J��m`�!�؊w�����k,���jCߘ�|�;[8L�P��˄�B��!g�>�Q725GÖ� �� Yt3C��}h߮��E�il�׻�f�����)��y�G���R)��� ��F��l[b�4���{lp�~ û�._3f�]��[�L"�E�IE�\�e�#k�c��N�ޱq!�ե�;���S:5���HZm�'P�#�k�� L!�5�]���62Wo�ŏ�T`��;��8]�0;�]�&�@;s��[^���X��j¯�B�<��#�0�qҹO(46;�}��6�
}�3����������m��F�h�Z��o�\�o�$�3�8������j�J$�F�3�̄5�Hpl�|��@�\gi��ߔ���k��[F��R�g ����x�=�"{y6���%��`�$�2�� ��цe\�O��7N5NUm�' =3��+����`�t4I��Hˏm�e��o�d~[1�]��a�i�1�m]�,��sH���M�H�D/��P�� ��R�\���!����9�}@8a��ё��F-ރ8��X}u$��W��.��g�r�%(��*���Pr6`tߍ��%7+3Q�D�jԬ�M��͞x�����
���Y�`ƅ�x�f�r�V7Q��yW������ ��߻v��ӫm8�ŀmk`�ꪈ�L�V�ߊ�TQ�D����d���r?#�k�GKX���8�T=J�}B�|/�&2W�6wY���Pa�ߣl���[aX[CX�z��K�90GuU��9����!�hƩu�"��W1��t��Y�J^b� ��,��|�r��OBn��3��_�m*��]'�h+�w*X*�wys�hʾԎ��N�j�ݜ�
��i�������?-��!�\�<o�=��*J9�@�|�t�ڥ"�?��PY���E)#���?��N��B��.�I�y���:O�3�&>o[2�5�?RƬ�I��&
->�y���G!�ŷ����{�:>/niO���s�)�C��Q`����\C���>q=-o�m�M�a��pn�0vf?p�Q��*����<�%�� N��"DGr�N�eP=h{IZ��o�HE�S�#P�B�	T�L��l��ꠘJb��_3�ぎV=H���m#Ɓ�U��v�jH�Y,y2Q�*��Ԕ>��Ef��%ݶ����`&$P��}����O�ff�������k�3v*�B!�U�5~%�'p�XUҭ �"6���������g�kt���x��ԩ�AS�H�Yk���$`�\)\bF�s�H��%I�� �S��DGj�p��A��~d{H�>���l�z>ZxcݵOzN�e梲�6��*��qA�X���άO�s�Ѥ13� (L9~��c:����iU���Rm(�^�f�n�~\�H���E��/�ރ ��h�<��� N�[;i�:��!o��X9]D��M�����{ɶ\���岙��Ҏ�l��@�Z\�RP�j3zӿɆ�b)�M3������u��������'����Vok�R��)W�S7�Q�/=0�%�,���f>&������)���OR�q����N+��gT�4����N�:�	�����@(ٸd6UY
~���/�7?�$K�z���27��MlâO]Y�V���H�~�|&!;@��z�;r��<�Uu��.ne3���T����$���Xa�
�z�pJ82=�l���Ih��1�8yf*`(0�w5��u_��rH�r��,�A��
��Sl�'놋/���EG�?�;MD����G�(d��ꨋ��q���]��#�t��c��������^�*�x6��m����D��U�Nr�z@=wP:i]D��D�f�y)zf�A�.����QJ�W�������y���z"B�Z����1�O��mgK���C�V��L��b�P�l�R81�L���ć��ӁAI�������B��'	�Ѱ��G/GfԎ|P��P'E_��19����,�X�8�eO0e&� '?�����Q])v������(��M��
�q�Q,7�[g���-}���ݪR�D�4�G�7���~�%���l!�EJ$�.
���Y��P��� ���AY�
a����m#.l�ԙ��&��ފ $=%�Y��A��{߅��+�0a�Y3a�>��xѩZ��9Py�2��I���Q(��S��*!_ؚg�}��7�%BjI7��G:!���D�#U⥓��8�NQ��L��+e+��w��#1qD|,�����Hg$:�� b���fYx��"&&�3������Fȥ}��_$ݛϤPr�J��&����k,[1�$O��S�"�y��Ƿ���ߌ���Ӆ��s?N?�\GȠBy�S8�������Q����_�R#2M�S�L4�ާ���N������ۄ���l=���Zݸ<Rl��g�f׬yT.�(�֗��,�ލ\7�Sߢs�aIκ��t_�	�����<�e��K��܏�������%���/����U��X9
�I�g�e��P�����o��8��(j]��t�e�◨��ǘ6v/
'*���`6};!?!�ъ�Cݎyɡ�y��n�V]D1~�$�����nʎ٬��><7�0���W�C�>0��"��k�I� }cFR/v�T_��f�t_�y��M�:�7�pe�Y�:m�UB��Lڕ�E��ɽ������I�t�
İ�7x����r_fTT�8k��3ӈ���m�&Y�&��F��!!H~񻴊R���Cլٴ>�í�zYv,�;���z��}A�������6Ӡf|��X���`~1m�4��:���}f~I(G�o�d`��i2)t96�����]�U�{e�e�M���L&m\NY��9�,��/�ͷQ��f��	_�����ZK�H�����ñ�^�L�k_y���gG�ڱmXZ���~���ryƏ�3�U�P��*t�A��W�m�	�!��Yr���
����3�^I�q�ܑ��2V��x�}���V��W���b�����G��,��c�<�@���+мeC���%r����n��;fc�Y��bl�RS�E51`������#�\<=����}�.�f���d�������t���ڸ�y��!B[]ӥ�<[m�@�	WQ�'�h���8�{˄��u,�W�[��od���F�4O�Q�lNq��1WhX�21[u���,T��ͳC�/��ZE^i����N8�-��>�~�"���4����d�i�,6U��T��V�88�̿��QA�9R5� z���#��n��oZ>������9�?���㏹���gi��onƟ�v�1V�B��v&k�ݬ���2|΢�I7��N��l��R����|*7�pq�'���[<91���:�E��˵�X9�#��j�Ϧ�������#ђC8���38q�-�`�[�_c�͜r@���5d��zo��3����Kg�-T!h�
C�.�y��-2��t)���9i��B��l����w�8����Q�,����s+���@C0$�zD�l�7�%����3�L$��o��\��u�`�w���>���禪L�m�+��ž+�[{jzv�a�N�|3.��>?[!	�5tMg�]�Vy�7���l d-^
��.́*��V}�����$ʌdW5'Z���ɼ����>:����MQ�T���|F����{Do������t�u��נ�θ�Pgt!�7�7�u�:;ךF��ڼ��<�L��c
JM ��Y3D�P(��*b>w)HU]��~墽�Ƴ���4��Wz�p�����8��}�a���}�`� Vt��M��G0У�g���*2��5�l2'������6�v�g�+(��b�tK��Μ\�7���B\F+��Q�΅��o����`�B�Փ����1q?Q��Oe_>���KkRF͈u�&&�@�Q�K/s������F[�j��E+�̻�ʚ^���ǧ�E��}�ϼ��ۨ8 �)R�.��[a��9
7���K���k�5����թ��.N��y_�Z��y�D����0E�����	�~ɩ5�I��%bLo�J���џ���������.�y�=M��TH���->Z�m�gyl�,CZ(��#k���NhRs('�lRIʂu�%�KR�{�́^tK(�����%f��=+P�5��a�5�6�vKT�#���- D��7^�Ϙ��1m^�,k��T, �|Yu���g����ֵ�������ƤR���A�e��T�����g��u�aT������1yA|h�"�x�5O͉@�u�$�9�m�$+b�x���ϝ��ӛ�!?jy>��A?'#�}y����曨5�5|,�)]���O�]�C����7���:Ky�T��B/�d�]�-��Θ\;����F��72?�=>R�u�t�`����� Dڃ�m��Ƹ*�ѱ�_K)��-;�fާF�nL�xEp?�|K��h�4TF<R�<���n8p6Y��0e�"	�Xnx�N?%��G�i6���yA�tLtq�rٿ@S.�� �|~)S�>�_E��m�W�>�H�o5��m�JO���@�HU?n/�!�^�>w�����7?;�]�F��h�i�����ǆv��l��j���Nn��>~�gAG"܎^S5�,��2@sN�����@�z���=���5C�Һ<4IMsG\X# }tת�A%���0RL޲~Xm�7TLQ��9���Փ	�g?����C��SK�*:o�B}4Z��9ϡ�?A������fpj?�U(�r�(�랓y�����E�5ׂ�#]Ks��/$wj��C�!�b�xS~�	 .`���¬H��:���{\%GcxG,P��nd�N�W�ـW�$��\�#�2��{D���/�X�sE��f�>�+ה�G��D �`�����)��R*@e�k;|o�2pZ�y.h ��ő�|.��1�?�r��l���>�,�d$Ԝ�z
�:�Q���~�-6,ׄ�*n1M�vbm�9V�d�D~��yeB���w�LI������n�8�L�L�Q4���5�w�o��n9-_��]��W�Ľ����C���Z�GN3�$��k�I� &�<�m�"���b�q@,L(�����.k�m���Q�Ll;������������dAK�\���e��h�i���>����ћ��~�G�.O�u�kt���j�␼��`�ǽպ��
�>e��Y�Zփ�Q�O�B�T�B�J��*�1�Â�P�C^ת�I�z����92U�Mh�`Tc��0h�E1H�c���

~exG��"3�� �������4��9�Fg���i���Z������MVާ���j8���B����:�
�-���X[�NYi�$h��o�69(?���_����&���u����5�Q�=�e����E�����u1��_��̊ԋ��A��j�"�3NL����
�Ћ�븏���	�"�C13�Y�'�lAac�Ջ��V�*�����gy���m���b\�3������	�#�;ڹ�w�;�z��Rs���.���>�����	Fri�:B�χ=N��=�,Ɍ��~�	4�}0Ce#]�HVOSEsYv�y��ʇ��-M��0�?I���&�T�S�\6A9���8�}�Z(��ǉ�l�*Wԉ|6 ��j�����jO��A�+/��Qc�quF���Fh(��.��s�/R�^+�${nJ��M� �]i}�u�1A����Ul��?��к�Y;
�@�y̶c+g��t��0����hDw�7.�����,w_Z�Q�|�1�{� ��îZ��K?�Ϛ���,8ˊ�h{���W�R?r&%R��D�U�%�ߔ�����u��	St��$wB�%��R*y>����Pg����`��D�`� �4��g����_��t��(� �0��c�xv2 ?!���@���\`3�Z">�	��{���헋v���Z�jh�x��C�ƱDU\�Pf����q&J܏��}�g���9e@@bl���j)U9趞>�O�a�E����|�l��j�W�'?a�o"('�{�����J��'��@���Ⅺ+٤��0DI�j)Mc>Q�S�#�.�y{�kF^!I��5����"fLJ�<�4dC~������uw� $+��˽8FӔH��?51MQ�f�k�(�;�c�`�iF��Y��ʻ�����:���S�ԋ��)VжF��D:�q.6���"`�Ǖ;a�-�lh~ϡ��3p��.�@6dB��u�t3���\V�yT��;@��F���w��v5��o�W!J܄rᆿ��v�c���Ot��M�?��mt/�o����/�s��f�[P�%��j�xd��:�t�����v^o2�|�����ċZ�t�d��7 �j($�?�+��ˣΔY����G �)�������(哔̌��=N��H�#{x�3J��,�lh�L���Q��+)��J;3��{o7Z�(h97\Q�(o��4��1��鏏�q�,j�E|�*��9��Y��{��7T���.IK�	**"P�A_(Rk1�?���'H�H���	>|�P��c�2A��D���ޤ�,G:���k�Q6X!@�N��D]wyϰ�H�=����m�h����w�Β43��5�����f�CA��\��v��]��
�!V�*�y��㐽��q�@x��[� �+�?�jy&���.9Xhu數Y'6~Sqݲ��[.eT���sv� �#�+���u����A~R$w�3��Iv��O=!R}��!#���߁���!��L�(u��]v��
��M����hB�R�h���(�V�Č��y6�W�y|'4�^��IgAxܯIQO�:��ȥM�I��_�|���:,�bJ7dSZ�9�B��
F5Ty�� �c�����a(�o��I;v����nǰ,�q�|��/�(��G�tx~z��?���:O�O���W�~��z�y�H'"ջv�r�SW����KHtSX�r)��S���[��������$�H�^龤Vr�3w���%/��h�."ԝ���פ�0�w�t�ڤX�����UL��Ys����ހoBTPY��B]�B%�RJq�S����`���
��Q����d��ʝP�Ӣ�n�����_� �A�wh#\"��z<	�B�lGm�,��3�r�-�����	lya������1�'�PO!���f`�j<Z��f<���	qJ�*io=y�h�;�c򇁣ךz<��x��Q)�r�����[%*�K��aZ�~I�4����}[g��+�N�"j�9�҃���,'v ��c!��$گ�8jQ��[gj2 ��+�=�lwrA�b�)n����^��5.Aom��SJlZ�V{@}g�W5���M�\~�_1���f95o�AREV��]�0���p�ά��)!�g'��%:`D�V��1$c~���7S��.�.�o�������ym�9��x6N	
��<�Sm,)�T�<gfQ�ְ�ҡsg��^4^g��U�o��&[z�>�IB����rJһw��<}.5�� 3�p�G����^S"/�ʀ`� r��NHҨ�x{��Q�vb@�DN�Ŭ�&ex�	���<�������و�78ټ,���G����'�)���8f�Q)]Mԟ@�Q�0�inh���7^���y	1��$ لC�0����t�S�ɶ�c�+�Pa=i�v�Tz�r���IA���xe�i��3��A=��]���M։��z> ����Bt�&�]jODA�|�b�#��{�MρG�z�1��
~��P�Qyt#����s���1y<4�xBC���"���q�?Y��S�S�X"@�r
S��p�=o>[�eqY�jV!B�U��d/�A�pDf'ۋ}G�0�oPbB�4�D|*�5���H��*���dZ�&����DM7�Ho"2�p�5d�g<�t��򪆑�Wχ/>׍���"˖���b����p	L�V���q�ŸP�gӂɚm7�ƹ��s�`?8���k�iw�N�������`��SL���:)SX���K���G)�}P?O+�=��B�7�0�[ڕ6+�suvŽq��,�n-5;�HjX��嬵f�Ef���z�������{��d�C�����n�m����1��v�P}�G"I��*�R�T�L<���L�}t��ftT'�GJ~OL��'����ᘙ{�pqcGh�D{N�/�ą�P3��;l���a��7t�����A`�nkO( jxS{im"�`�!�Uc1S��\|-��r�`�����j@i����!dS�S�QF��.�mޘ��~>�b���&cj� ��\��V�d����X?1�x|ȕ��.K���֡�a����J�	:�x܊d���Z�d����+m�uO[�vz���^��� b9-�#�/e�-�A[Bʂ��а�8+�Р<`&G�����F����n�UD��i���&�(����ߘ��FZ}�BS4Kh��r ��󿸫�ӹ6�_I拜t�������x�+����J����[�`��}f�m�3ťv�dǳ�:�=EɛfLP�i>�'v�ܛ�Ԋ�7+AN��r��|�Lc�S��P�:��>З7�v;�� �j@���X]�j�tkT�w3�Z`rvة�t�@���D@����k>�у\�O̪#HTx�ߑ6��p��X�*���&�6;LGt��;'N��mD�Q�,�L}<�씺��B+|�G�i��t��ݟ�����ٶ{]x�[���2^��bZ:=�����Z*F$�Mq@����@�']%�kx����2�t��V���^c��(j��@Q��"���Km��;�J~�|Tr�4R�1d �z�=����>�~�$
3]�[��[[q���li�&��>xFqB#��!�T\��4�j�G�:d�ħ����А�����Ec�T?fb;�
xa�E��P��3r\t]/���%FP��PV�k�Z�ۙ��H8�a��xW�W��:��@;ұ���	"����߇������z� '�j�Ƈ��W����bʥ�~�F��`A7�.���m{^�_ssʐ9:G��uԮ�3K������6��5K3D��*)�����]_�ϫ"7g);�z�>υ�[�ɐ��.V��c����Օ�g^r�}>��\�u��"z��'lga�g���s�w6A$h$�3CR�.)J����4N��o��kn�a���o�*�;��@�''�'y���A�+݌PG�+=MDl<�ܷ2��>�8��B���Q��÷��R���w=c�n��oD	�~���^��{�@B��f��4Nz\^�0��C���MC��D��~@\�õ�XN !����5�\��� �P/ڰ\dz�OKL���D[0��*�YF�C�a��{ۉ�u n��y �3q����R%
�Y�tG��ïY�G�t2Ϻ�u���
�8�*Q��ә����]������nѪ���V�	6�\ی�����JP�je����`���;ĆW#��i��*Zo�(0��ܼ�IS��>CCo@��*���0y��N(lcL���?�>��l�+n�|��Yʏ�h���!���0���dbj�I���G�2�e�����(0]n�mK�%Y-*B��k�3ꠙ"	�a^�x���).�j0=~��i�\�����͢��'�3�X���Ā�)o=�v�U���i���e޼V�� ��� �O��VgAj�x�#e��4gw��ʅo�R��4r�Vb,��K>'zFd3��U����2R~�c���0�_Sg���H�'~�(X��}y�Uw��Ykg>��WM �	P8 d�^����.��g��k�1������
>W�b�a b6:%���_�/�j]8	?Ü���R\'�pu60#̣q-�(�����J6R1����4hH9�ܘ9\��7֛�-�%i"�\����q�~����Hһ����d�����ű!��\0w7���l5z���BXnXD��*��"��*��U�F���!H�(g���-/��f`�5VI'�C�V��4����Q�q>mS�k=�4�m�=�Z�H��$��'�8=�d_�-`'�NAf0���㭄!ཡa�'w��)EH;�I+e.6�#��N�gz���$ן�㷋� �.�(�j^	�\����?+�s�7��
����4ak�J��i�CX�|����:[J>/!��-����y"��$JQ�+DB�����n�)���u�&���01�N�m琢��jj�
�&�{��D����֜/>�AØM�6��M�?i[��̵{ �>����a����%?�;8	����&X�����D�F��?A���3"�a��QfOҗ�ꪚ0��/�o�p]�Oi�����!1}ҏ�����z�����c��tsǷK��yR�,rn�i�D��?�e�鳄X��Tb6�q�xߵ�R�A�j�mC�o��VE8�S%���j.�
[�a�ys�*�䃝�uˢ`3�����@�g9�e��ķ,zȋC���=�[��Ѫ�����5�����^i��\V�;��΄Y��.��9$(���j���f��)�hdCC�Lp��^q�%셊u΋Ԕ�'�m���������b�ZN�ZK:V�Z��懠��E��q 6cm5:����o���Z�a$��` ��������V�d�pd��UHƩp>!%-(��g.�̟2�0�C)������ףZ[��<_d��p�?�ء޼�Gq]�ʨO,���:u:��'�oȤU�"wz��6����[��%�A9�ޱ5�c
�� ���1WH�_�0-���NΥ�#D�����f�����^����Qp�`��e�f}WGEo:_y�7u\]0o�-u�P��>�
�³Bþ�S�<{n�U���6�~l��h�}ᡓ�j�����I���]�0uu�\fd�Ez�@8/����%�3y����aZI ��"k�L��D4nt�V�.��|�h�����c�'�?�[ ��7��~͂�ӿ@�m���mR� В�ؙBЛ;�5��Hp������W�e��a��YU��� T��Nd�e���Z'gP���M�c����f�zb�];�句X]�JQ����ݵs(�U�cl{�=�A��&j�u��� (I1X��^nG��V
�8�������,2p�xe��<�i|F�O6��{c&\B��;�V�b������h��D�Ix�����q�|ؑ��Ӓ}_�0�^�.ͫ�pB4b����)(S���5�;��b���%����F`����0����g�9�P=��WJ���ƩB���!h3,G��YM}$ ���/�,����Ie���6��S%�J��I�܎�Y�1k��C����A�>XA�����g�H����G����s���z>�Ā�����?���k�b�!o��6d�=�`�U�d�.i��O�,�;H
�$�M���x���K��J|S�T��G2�i���=�,��t����{ʈ��$觌�׏�F�(��꾲��e�Y�X��<�����E��/�����)�
���r�۹'�r��Ol.DX�<��0р&��9or��Y���k�@�U�œKi�����L⒡JH����W�H����w������΂�,Қ-Z-���kx[^k���B�e"μ+�v!9�'Pd�Ίa�/M.-e�H$@���?���z��fN���Pq5�������-&��7�U�x_�E���XZ�kK;��ʆ�,Z������_O�5��3�\���}�����HI��.���q�Z�I�����h��������-�_&0}ODk^5�c��	z���H�ÐB���HWحe�E8�d��͡�!�#cS�^ n��� .^c���]+�95:$���,��� �(F=��X<���m%QC7���4(��xm�H�Ԋ�3���)�n_m�Eyb[f?�$�|G��5��R�u��Q�D�f��<a'�Nh�h��5���6	3��u�Fm�n�$�IQ'l��0�n'Z���Q@�C�w�_  3�S��2�I6��z��Cz.��l�z	�I"e�ɒ˅-��X���N���	z�v��C6I�Bwb�s;��-���A�1i���Ġ/S��}w�u�Ł1n�@�7�ykKR}��>�,��1� /��I,����;ĠtA�i�ݯ�r����(O�p�P��3�����IJ{j������)8�a�5���t��h����Y�jx>\��yg�Bi�b���N��F������)s�X�9�Sg�$�0M�]���b=U�H�r���e|S���ҫ�U]F��0�|&�R`R�L��٣�V���3��J�މj�2����=@�VĤ��2_�@�y�GQ �n�CB߳�\�~��ˁ���S��7|��,�'zes�1�]��\OO����:hM�X�g�(6i��#𒑢��Ќ]�zNw��2C`Ŝ2�=��R��H��s�ߞy�w�_��z�A"��~/�!b@�b������s�&(�jˉ�Y�,�S��ǙǛK��N���ohP��@�1�A$W�2��d�ĮKy�0����i�)NnRNɵ2�@��{��$w/|E0�-��L�Q%4}mC�>�D�T1�GuG���Z�~6����x�s�_]A	�>���C>ئ�(H�Q�ǂ����u��c��b���[J�,��ױ��G������|x������V��-!��F��~�k�f8��$hP�H����s�� � odw�b�Ga�y"�E�4މ�I`iR�1{7�7O��8�L����
X�����$o�TGRޕ�mx��m��~}�H�0w������70#
+�:Z��NH)� ���<���].��PB®<v��$S�������T�~0f��+gVT@���A*L��T���|W�Kh�-j#Қi�΃5�Ѥ~�G������-�ra,}Ul|ى��QwA��7d�̈́Pz��Wz���;(�ɡ��/9��J��K�Xb`3"�)3V�oڋl�Yx��)�Kz�*�$�~��<����9�m�(����}k=ǗK⬘l}��TF�,LTf�2�-;Xe�Q���<����doIv�j��1���EY�2�B'�b�Zu=����K�����9HP:���B�f\��X���"��W�i��-xxc�Ce5-$�7'��A�����
�#օ�*,+��o�%36oi�ē�������rCNO�4�����I���&F|`�'��w#+c��W�͓R���x!�#KsM��U�wp����5	�E{��7|׻@���z�Nx=}�A���L�챴�����A��h�۝kP�l�umF"�η6�y��[h��_��5�}�X��D�vc���>Bf�.�1��0y�b�@љj09�����w�G��҃��$%��) >s³(�wt\��h԰[���J�"ǲUQ0֛3���6�k}V�\B^�M�����t��cc\���ȡ��9�j4�٠�J������K7�S��e�/��%5�&c��inn��'}3u���*�9���[F�d
>|�/*K�yO1�]�{*���na�E���]�D����UB� k�F.=��?id��d����3th�ȒnL ��WH3z6a`z�PQON����,�p���R�~4Gb7�U9H�Q�������M"��@�`�Z~�7�)A)�DP������b����p���u�4' ��E�D�^�緯j�hr��Ou��]�\f�!������S	�^�\�J�������0�,�9����|L��gN��W�ʸ�%o	0�r�p�,	��Ka#F�Y��	�Ч/�M�p�Lu��Ց�'�_'�|���
�Ǳ2D�%��F���r̄�ڳ%�=]�"����6'��Ke�d?IE_Ld]^�i���\�h�3"���(ؑ��]����9���#�5p�1m�H��	�ݎޙi�2�'�VS|�^���C73'#��!Y���,Qr6��`6��6X.�-��h��'�_�������k�l�J��AC9�`����ҍ/�\7�V�4�J�clh��l��^,Y������Qq���C�L1[n�,�ޅ	�dT�����,���|��e E��=ty�ɛ��(�i�瑒��"�>�������o�ߖܻ��B~�V�&#�4ߟ{"����F��}c��ȹ��M.���tri�G�]����@��v�U
���}
s/,.�0���^�q�����Ks>�#le<1���������F���տ!�P�m�D��QcL$Sf�` E��qxt��Y�Q�����Q�\��N+� ���i'�d���u��M�0,��2?�Nװ�}�9�v��!j7p�y�A#�+yzXc�e2y?����=� ^�'�X��=��(�ܖ�J��g�	�2��.Q���2�3�L��c��dz�-jI�����C"!���%\��=�Wt�vh����%�{�S�ͤ�t1ۭ1�
�@�d���B\ُ_,ᦝJ���H@���4T�� &�M��ؤP������1VYkQ�
��Itj��dZ��~��2d����EE^�=�rG��_����Hܰ�.���]�]�G�Ӎ�T�{�Zd���b�L�����)����K07����s�4�y�S|��*�}H�oe�\��
ubO�����xIc��,�~�"\����3��9nͨO�_tڀ�u�Y�0P�j��ݲV�]�w�G+�
��iYT�t'�f�IV�bp�3(Wn���(�6I�פp�����<��u#7xVY��^�>MExA�3�o����uš��xF�� �P��.��w>��k!֙ͺ���#D�S��e�D�[���O��U�Jb���
!�����^L�S5]���&�l�p��	@�N�˨�;oU��#�a�N3N���4qZ'�`�R�}�K���e��x씪����F����_��^T��Im;� �eZ���HH?�n�K������� ƚ��4�k猦X$G>tA��'jp�ή~�W�f�/:_�BOS*���V��B��/��o���Z�'`L�[��M�y�P�cP�D���G���z�T��v�$�~v�~�U�e�d�%�"��j�Q�@����.i`�g\��m:.��߭����.�M}��+!)��j��K7�4,�\s&�h�`У��K�s���=�|XNk �}ϊ-ao�-W"S4���s�"'R��c�w�����Q����Q�ƄbX����78u�O黲� �$ݛ��~˰�	��]�����W�Jɱ��7a\v�pĲ�)hr�OGbb�����@���(��¦��cftr������i$�솭��U'�9�X��=�h)���D.1iw�����d�5�vJS����W�����9����iA+�d�b���<�km��%C�b8�<�9�.�k�i��N��.�(�輡�ۡF�3r2��O�$�*���oI��VL��ς�5�}|�Ǥ�S ~�����~���G��6+�hʽ��.�Ӹ�ٜ �ǆ(�8�)' �=��]������ƨ \|��E������i�p�cb���D�
ܵ�Ho���2�� z�㉤��C��&�ɉ+f�V@-�Oz��\��$-�I]���S�a�H3/���$�P�O0S�U)�WȞ G��[1ҙ2��vC��Xt�4�W��]=c䉦��6Ӑ�;���@�oț,G�o�GJ?�Ejp�̛��/>A�Q���������ۻ�۶�S0��t<|�<$�}�$�&��5v�������f����u���E�F��e�T��q�a��M��<�)��Hib���l1�Y���QP�����
U*Of��XKZ���@hX��c�iHO��)y�b��+3AB�{��;�Ѽ���M�8����O�ccE<dZW���Q��?�?ؚ��瑠�� E�3Fӈ�8�˜@=!�v,��(ã��GWӐI���ى�W��Y_��dy��t����b�!�'k��>87��@B��~����b8(|t�����17�a4��O>��g_E��o���۰��5T_ߧ4�8DD9������p��BЮo�p}JU���!�7"H�o`�?�M�~��þ���-/)� K!��/��JT%�G����N��n�oD2]p3�f��L�_Ϙ�l�e�Ta�&K�#|��kk����p�W�A�h��T�7�r��v�Ec�'u���2���yI����S�e��G�\��f宿{���Q���h6�)��x�	n�ߚW;e5̌��y�pŻ����p��Q��-'�����|_�4�f}A��Ic��1��4��=�M��)����5ڱ�n�<F�?�l���&�_���T�yY����"�l��/̜�1I��6��d�>�!����E�*��0�%����fe��/����YNlV|0�P�N�4w��,5����t�|��Z�PQd�(�БQ�8&�xD��9���9���2yo���"0���}���� e[�'cib+?�����`��iǻ)�F����@U"�H��;��|a�	-iԩ�Mc�E}@z���N����qg�Ħ~m��#'��.�׊3)>�8y�;��9�\���v�^I�C4���������[�:��I��kM�>�gV��M�w4:�~���%��,p<��~U�$�_4�� u��yc��C��@>5����{���sИZ�M[�yFP�#5���z���
�G���B��½E��B-�}^�ə"DG<�%�4ꂂ�A.�n��i�1����g@;�0m6�Y9Xi-on��x�Oꊐ�֣-צ�P�:��	'�����D�U
�w����@6i���f�I.�!�hBXD�u��!'�~������7�p���|����cZ�20�i��yP���Rx(I������Ӽ���%;�k�:H��8��#��W��x��b`7]�t��3_e{�/ ku(��B�<�u>�k
l;b���ˏ�I�ݎ��u�6�QV���QT梞8�j2a&4�t`ӗ���rV��04W&�?;�V�b�;`�A9ղ!�|#o<�Y�)��~ϊ����[T���f��_��9��"�n�ؤ~���i�7<��&'�3����!��
�/�ce�'�c�@r��	��)��20av2_5LR��K`����^�I٫_9�ҿ��Xp�/x.�]Zs����o��ՉōRo��;D"�Y�$��?vR��1�z��zepM��Ό���(�	Se�/�sAɢ�Z���/?ߖ��*L#O� ޲xd4�^��2Ta^�B�0�VdԽXe�g�w߾]�lSvc��|O�$%��gCw'�Q�z�ł�z�O�QK�nzU1Ҁ����1�2����*��axE�5:b�֤�
O��z��B*���8��t�&��� 參�@��ly_CH]�i�z�{.Ã��;y n�$}	(UB֫T��s������}�����|��}`�nw&�i�Y��T��j��qJ�*69vgXum��'g�h)k�a?��� ����(`j}O$	�|�;��c+W�!�:��!�Ufb{�Κ,Ǔ桱R�=()R-e�n�	D���"D�P������w�d�{N;"�h��+�$wXR�2���-�^C���<��$�fo��Z�g�5�|�񅌢 �[?����@����k���U��u��i���9�ݍ�&��p���3�T��8~�_Z���+bLC��X�3l�
�~}?7�O`ı)c�a3��b���?gvr��✂J�J���V�GRj�Ж$f�MR��)�{�X�dG��b\0t���z��!Zt#`h�p�����#�@�X�]�+�����?������S��d`�B�;q?�Վy8:����ڥؗw������0ǝ�:1woݜW�����1�� M�0U� ڧ_�!��ϗ�=��qhY(A�y1������}7��r���n� ��Y*�N�h�b��su�L,1�(5K��ܱ~���-]i�ZkWgِZ
�Q�����KY�x�*�������WK��JE3}|���M\��\D�tG<���=nIx8��XSi�U�`��y��[�|GR�7Tв�w:6��6��}Ǣ�y�i�����-���,�׹Ù)G/�)-2ƅ�TWFY}�c�=��!&{���.m�χ�!��5 �H�����ݖf:y����:���?�1m�IvR=�u�ƶ�=E*3>���h�\��:�9��-�W�\����v^8�[k�,��_�����&?`L�����e��
L�Gt1��m��[�@�v?����4��w�
Mv����R*�h�OlC'���k�`<������6�S6i\�ʡ9�$�\��x�Ą��_�f��z�f[��X�{8�
a} Hk���[gLB���D�O����9w�| �������?@B+��G��.[!_nPM�֏]jl�����5~ͧ*4��aVHG:ֻ��40��yd/�Kq��U�J�)l�P��Y�
I�U�����b��SF|�v�[�q
�yt�{<�(J�?'Y��!]P'�c<�w����v2�E9����˩��_��#�GO=lmG���K�|Ma�~��=�P��n���A�9��tTW�K�S����?�)�->����ӻc��O���n/+x���ϔ.����G��QoHV���փy\�J7��iY�E�ue��U�!�ɅL.��iM�n�;��>�\m�T�]��Uc��;��`g�@a�o7��O���� ~�?�>��E~�%�*�Ý
ݼ�Z��L䠦����rV6l���_�SU#���x��O]sR49�i�x('��-�;J���A��K���H�L�����m�y�?��f�7 {S�m
��Ņ�	�T���f5�������|�N	iKX4�v����|{���L1{-^M�|�A&?��禾��0��3QOM�R�m �6v@�O�
��������M���\4��K�]��`K�26�M�DVm藘�CzM0�p��{r89��)�6Q���R�Q�FU�N���Q��V��P���ص��|[Itu�n���P�[��|n��S��Xc\�.n���ГKj���r4��}l��L z�'��!�VV!�ˁ<���`id���G����e�mg��LU��@�*)����i�I�K�x�O&Ԛ�Ӧ^�H��
�Է1��$#I�`A-n<�u�S���+�_3rU��헾��R����[͉�5���bL���o?1�Q��������N��ʟ���������tE��$\���SV&3�g5��� >����5����!�
	Rb�D��f��>�&�m�.�tK��}d_L�ۗ�2�5<w�HN�?g���jJ�YW��S�wИY�/�
�|�m�D�,;��[�	�����&߾č-j���G�1��r])�ⱊ����	��bμ8�d���vV��G7d�\t����~	&��FqJ�?F)��A�0���.r�,<���e����sf~�A���H ��.bm#]�Z�浧��u���ٿۇE�$��'.u�E�èY~��5tkđ��a��H~�OBD������R��t^�2�?��.��X� ���k�Z(��bNp���|ў�N#r̀�b�k�������U�]��(P���u�ߟ_��UDp����/���IL��&P�I~
����:�����`eʅ��Τ'!,�o7���<��@��J�sīv�.h����R5�у�᱄��,g���a���Ā]/�rZ�<7�edjڑ9d�?��_qsfN��o��*��MY��z�#�]I�};}�l�w�/�ϗI ��m&�'��|����+4>~�tcF&��fG�R��w��C�ľvd��4����9�ԣ��_�5��Yw���r�Bd��K��S��z��"��=�[� ��&$�a|�?}S+K�o� �۾��irT,	����^T{ ��,����D�[��/���k-#���m�r�Hr1èO=��$<���7��Αo��y-gE�S5��>:2�e)R�ؾ��곒���}õC$�z����"��P�|՗�?���L��"�e��pvxbԉ�u���� ����!�����s���Ny��4U9'�8jl��*
-����}���`/�+	d�G�np:\�իmJ�<�*714��6�z�Wh�H��}�QN%E�Q��)�x2���\�Xx7ۡ���U��c?ȅ9�)L�ʗ�;��3jj?*vi�`(��S�Ü,��]i�I��Z�iְ�T��~�N!y
2�s�DdrB�[ok� 9���PE����	�\�j������-%���\^�CK=i)� Ɣ)�h) gԋ���_+�D�|�IM����^��#���I����fˁ��q>F�6H��E�ܜ���B�5H����g���b�ܟ4�s�m;a =�d0���%��P����!�8x�-�.M �qJ���;���xU�����J:�?W@�E:���_U��31�V�` 8ل:u�TB��j�����Z��60Juee����J�&E#�t��⠏�RП퉜�W2��!��E5�`�Gt�\|7��v1��&�"Ϋ�c���L7�.m�HH&)A�K��+ͦ(`��?-�ɼ���g'�v�P@�yֈ`��KOq��O�U�vj$!�j]�����u*_O4����C�z�~�V@�:4u����
�x:�/��v�Lj��v����&Z�G������C�����(L>wT����W E������e^�����`���9�4����F[;�?尡�A6
�9�h�j�����F�o|�~J�`�L��m�\�)pVU8�I^:���$�t2 MuC��
.s�ɞя �mg1���B�/��M]�cgF}M2��YS���QJ���K+@س�9	�ZUg�n�o"ж��Ǵ_�� �"�X�5xeћuKQ���M�8�`���Y�S��.~SYHؙ���ǄQ%$�g��A�ol���2���Z'���������4g��+����DfU�X`2��%�,��NJ
8��F�U��0�n�QGV	d���-���#˙~:��qL[@ٝH@%��(�i�2=e�-*qJ����l���6�(�\��������s�S���.FW��ǰ���V��m�	��0�9�����>�l����J���,lu�����U�.������g�4\�����L��$ �� lM�Za 6�Ӗ+�؛[� ��,\��%�6�M3w��#���8Z|���!SS�������V\�9�W�l}��$r�aؙ`dCP�,;N�bH?&1��U:^<���#��6�]�-w:cj�)� �:^S�f1�L��&��@�����e7*ٙڤ=�{<���
�E1��"���?��`�S�V �o�(�?�ve
�?<A�Y�2��
L�3����p�H��ꯃb��ٗ����/�U�;�O�G���>s7�Gq��K2�'#�fd�����a��Mk���e����� "��z���k"yZ��TF�R�m��_�AbS���g�%��� er�8 j��K��MH���P�Ê��N!cW�ޝi�GD1�l`��� y���,������!X�EQJ����a4!�lE�L�����jOd̐si�t����J(������	MpV�m��*��D�;�}W�=@ ���!_�[4IU��׮������E��A6�o����7�^�{��W�v�A����A���O)��/�����/��~5�V*���r`����� �c�9��\	����5�(�0��H�{��a^��<^A��3,5Xf�D�%�҄� � �n��`un�l�ر87C���o��9?-��>�5�~���Єy0���Z�=����b E��gN��� %S���%���w-IQ�*Zcrv��B��Z9���ټ4���o��W{S��;AY��C�W2��$�\}����T:3�\�B�
�U]ٻ�^5g�:Ia.-�3��r<�2@1�������S�χ��l�?F��D�d���W>Xm:�B)�b�O��ma��˱ډ���}{8�@�0��rXوe�� �*ZBe�2�@h���/v	t���N0$�Ac�z�E|7��}K۪z>v-ZB���䶦T�$]����,�+�k�)����e�0��D�$J�!ժQ��O�<U#�vv�Ov�!����){�Q��~{�Ib;|<����y	�<��s��]ï1'Û��O+���tG�����Wo��쥐�WLE�
2��N7���!�Rڵ�6�r��M���m<�h c۶O����=I鱣)�D+{��(�p��2��a����U�$��]�=�	z���h鳝 |<�]Z6x���3Q{� s��|������������>n�~_��h~��_Ճ�r�i���B�8J�?�)��dt7V(w�.�f�q}�O����K�2� ���N���lkdɌgx?[�����윾HRİplQe5�@K�\��[��� �<������̹k��*Q�N��ma����<VtgY� �!6>���A���K�;�� ����tG�]n�>�\�"m�߉�V�&p��� [Z�]�U�#�@E�K�It���}��ܰX��T���i�i�Q�_1�צ�~(���&��wq�H����f�'�A�t��x����pͽ���րXv�(�;,�"�x�����5�'C�DV�y�����3��p8�+���a������)���:��AI�u�w�`]�U*l 9#9���,�Oy<��T�a�8�K�_,���ߢ���~��s������AH|<�L(���*+�ȋ��O�O9�����k`A||WƧ��qc�9�!
A�].�m	���'^	T�UI���Z�����1l�Ws�p�8W��w�:�$�*h���溳}'��0�:��]˹���1r�,�嫰u����4z��sc%�X����Q
��i�b� 5 �RM�i���q[�_/��-\�	m�F��:%�C5R���Sn�;1d��]*�5d�wy�b:X](x��=�|��m��˔�5KH *T��n/��h׻�����y�5���Q[��L'��:и/����:�o��m&�CW\o�Y��\s6��l��b�@��J樂U�� >���@L�wΓ^��qQ2{i!.�\��	��X���.�<�l�,����>��6f����\�&���N��ö ���. �����T��x��N��/�C`����2�$	CM�(��7��L��o��#��#�qm��+�QZd=�񷛷�7@�X�wK��-v����K'٨���+�v �44��&mٷ+�`ۃb�� �U ����M��ǎ�X.鳏����Gm̽&v^��H��8�������_Ɩ~&�~�ϸ��0P��^��g]�0=?��%/�je�@�������r��=�O�(�׋J,��9nS��k��<�_	k�|���_W��
?�B��M�+�<���S4�̤��2Բ�q���t�'hP&�}o������L���U�1�+�t��<�R���P�d�D�sA�SA�Ȩˁ2�H�γ��RY!��w~�s����|[[�+��:*�]�JQ��������Yt
�9ؘ6���<��-^#��JC�o�.{��Ma'<%o1:ɸb�]W����q�@�� zd����g]��G��jo�A��=��6�=2}Y�����~��-���SH}��j$\w�����L�<�R���iH
5�ߨ�r�|~��cX>�_�I�·v2zgm;�*`�$�h�FH�b��pC渇�<	�t':����Z����'*x�QS����.:*&i�Un�T�1~�� ��߄ݭ�3;��Q�q�ˮuF�� ��D>�Vw��#c/��`glp��8�4;V�a
)�T1zAD�Ttj?C�w�����1�����/�8��;�UQ���]��u-�Py��bTY��������ˮ�qo>�W�p����$J��9�bD��4>]�A5 ;Z������S�ћYӱj[�.��*���Ȟ\��?S��&�4���q)�y
`����B�zhxU��'$��Ȝh�Ib�O~��\-6ޛ)������V�O�=?��_Şr�BC��1�c�%I�~�F�BQ���(��.�slT�/3��B�\�#R�E��X#%��x������B@8^k5��`d�� c@[�����!�&�(N�s{;j٣�,.����=<�j�\`�ӛ�
 �9�:�26�4bj8v�x��M�J�@����,&�wƚ!L�{�(%l0!Z��ݥ�ڎ���ω�4�	���묫�'m� �<Ʀ\�}!B&�7EBu�Y]��D��`y��2�m)y
S*^��ꢡ�EU��6V�dp6$�vx�qp�+��KZ�oU8���JE�*\>9l�|���T�L�'���*xz���KsV(�S�?VxϊM���2>�b��r��V�m��J�'��P��OPs9z��Y2��5V���S�����S��Vg!�!4+��iTc�]��H�HU��## *�mx0�B1|Jgu�N�xş�
泶��>ㅸK�)��{���̶��i�������X]w	������@�D���t��j�Ŏj�'�ڠ�F�o���m4��"��8F�kW�Ǣ�'��q���;������������dY]���Ib(�h�4˚T>��
���j?�;:@�����rX �jڂ�f�V� ���<
�fCY�a��t�m4��{�^�;f�R�ϴ��'qq���l�����t������}�м��Ą7�'8f,[9<��:}WX�.��Bd��)Q��R�|�`�7�� ����.r��ۼK��3�L���١��^1IZ�x�kl���̮mw��1���{�7�:��c���J5_���\�y��)��ك����#'/��j�����,��Gy��ov�f�����ب/K���d$���'�m��1>l\���ŭ����KY���5�L��{��\�,.����d��a�(̅jH��rb��|aހk�T�N����{�؏��q���� �S�<S�- �2W�C�I|�Qw��u��t�ش��
�	 ��/q�Y}G9迻e����@��B�0��L_a�
d�Ъ��Y�kԠ��E�q����~�~@�dO�F�"
e�e"��q����w�h�X�Ƽ�UԯB�7�4	��� �{�`��5���H(����@���+8��평g=Ya� ���s�5�A�S'��4���G��k b� ����~��p[����J>�!K4~��|�0��U�Fe^J Q�6T��O�ǥ۸�g24YK[��|�N��j�k�Q9�h�pO�g��֒eu�sa�<� -$�}�m�/58��.����R6������d����ߩ�T�Y83��[3�-��p��a�Dim������sP�N$��v���<&6�SNn�Bߓ뙧�n4�U�0��M���h��KC���\wRxD��e�	zLQ�#�Ē������t�^����)78ܩ�������S�`l08L�	Y[�8>��$�Ͱ�h<+��Z�a�4�5'_ b�R8����x���IxrL��64�&���D���j��Ht��R9%�:�R�a�΄��94~��v/
@��4�S�G����X���%���>~��f��h��"}��AF�s#>�c��Gdr׈����-d��KP��6����ℿ�p��S���4-0�H���6�� ��]��e����I
�ߟ�l?�ై��]n^_@��֠��R�pz����_-׎��*w#��:zu��y��ۊ��d��2MA�#-��휊��u�����4��!�o���[j�^�|xPԨ��?[֊���bGV!�p��An^�aC�#t��40���D������*31 �ݲR� ��������̀;�n䖩",��ٓ�\�P��^ ��'�T���A�TA���Ɨ�����`�	�X������W�+4��)L����P^�w��� �x &��Ǟ�)�c[-RM��
]y�W�c�_���p`�״h�0_F<D,��{�ek�K�J�@8mZ2��/��~���ۜ ���(-�t���Ffɉv�5�p+}�P��!BZ��W&�Ҿ㟂��'�w��dO��/��$��X�tU��1��_�5����
p�l/��Vw�+�;�:���oE��G�N�\�r0�h�#�72�J&ؼARD�fV�bs�/�Ľ WS���+��|6ҼռL�1	I_����}�W�,V���
�+�E:'<�(�1��	v�� �r�����J�� ��h!ΐ[!���C_�yl���}�-�%S!�Ӣ�m|�t�e�Q�����8,�<��숀m�g�~�,6�����|�/�B��Z@H%n��݌N��o�W�&X���F��Y(�/�BΟy֝�C��/yK��lZP������L�3N�R�-Xg2����5A�T��4��%C�1�D�{�����@�<�C�����u�_~e����R�f�Ip��M��K]�������/g_ݠ;�����j�`b�yYM��QĬ~UW;k"��1 �Cān��vK�}� �ܤUP"��^F�UC�@�*Luӊ��(`FࠧJ+0vB׹p�� PJ|{lIt�tN�e|v�`Z�NPBJ��0�K�_a�z+���.e��t���nh�����Ur?�gx�N�)����Ɓ�UZZ!�݄%�o�K�Jz�H�@�����Ă�֝�x�;�P_ Q�'B�ƥZk���!�{"y_ç(��a󧅙�2 ڒ���\��Ɲ):�&�'��}��N5%�aE[I$"}��]<�`�A�S�܎٫�F���ו�i7��X�x^�
��·����Qfc��$�C�o}�g�^da3ҭ���ҟPo�s���ͻ�e��'�U�#_m�&BsA7/wk��!;8s��睱U	±��<�����6��tX*�����fc��Үgғ�O1��U��^m{��I��כ��e"Ϯ��|�c!q*��'�R���Mx`L˭�3��������75�1җI�J�����{H'�.����@e�,$��Ȝ��,C������+!��Y�G�Yٿ-Ҷ��f�4�S��!�,�]|ϭG��4�Z��C�hE^5,-W�rlK��>�8��3ӄ����O�$��yh^�2���h�t�k6��#�5�>�p�{!���蓽
����͙�7���GƎ�^�$ĭ��z$��R�V�D@��O.�>'+�>xq��&>��h��8�n���$\�_�M�O��,��p�8�����CyLN@��=jYy��o��\i#I�a?�9Ǌ'"Σ������hλO�
���������:d!�ɽ�ZB Y�uH0Z9�%���,x~�5�p�W�ƪ��]v'�s&W��8+�1��w��hS�=Y�:�q�
.O��W�b	�CJ��;j���1FI������A}Q1��A�ʠ�J@E/_�i���Hن�L�n({~������w�CA<{�E��go.��%|:���M=�����>� �®s]�ȥգů��m똮��Zg�툥�R�ә0�ჭ��+/!���/*�Ui�Ţ?º����tyާ��W^��ˆ�xw)�J7���K
�ۣ���w��7Pok3f㙡m���<��ѳ�c	��V��I�M�׼];��Be@��J�o�$Ӣ<GW�"�����Vca�
�vPj��_��ru��� QgYsp����%(�&�y0m�:"��`��kս�6^�1�Hwb�j�Sm��f	��˘2L���R��h�-�knbyk\����y�K`���Ec�KT˪��vF������[���;7��>J����P�F2���׌��xz�g�n�Ł�
�m��8���w2u]�+[(�Φ�e}Qޛ��������9�)x/68貤��/>R��������QEЀ
۪�
�7�/WyZ��ؼ�[XQems��M���x"�5����)m�0�(���1�&d�S�?~�f94x~ b�r�eR�-`�^zP\�[�zjY�UB�=&�m��ϟ"s�xI�߬r�/�yC����m���DYu�0������."L^S p/SO��Vp�5ع�x�G�.�	o��T��O�
ތ�aL��7j�o����IM7�0<�����_���o��t'q%3'�0�8Eb��U�u�02X�!V��b?uю�j���l�!JL�r���0'��
��I�d�����_��yn�K矉=]��"Q0�k5�ᙛo��&ٯUf�b�:��|�-a��#���7�I��@տ��f�["�V�ic-�7���F�a%��J�Q
ׇ���'k�4"fRA�vZc{�u9��P�4J[���8����E8�}��OS��@I�t�� �ᗫ�*���
~��j�����	��ͣ�b	gH�����P������b
V��%(/�y���&R��0�U?�`2#�2B�>+�f�Jb*=T�CیMv"�/�����W��G͗��uћ���u=»��]���_���I$��n6�4T�mp/Y��5+��'��8I���zԘ�]�Fo�c&�[6�	u�/ܜ�,�~�'�� U٦�,<+C��$O�v<>pݦ�"�@�֊s����%]��Ft�$�dl62��,s�w�{���VC�q�r��&�zA9l[��K�g�7*�5A�4���r`�L<�x�B�W�����[�	�ځ�� �T��T6�M/��Uc�r���	���x��ƻ�8�wW�Z�)U�ە�Zd�Ż�g���E�/�/��y�<���<�����;�+?������o��H�V��'^s�D^l�¨��`9�[mp'=�ʔ��/��(d:�C��B�C6��jJb$�6-;�|�E��f6��;�i��>�F�[.���y�A�e��w�w��s ̌;����8n_���]7c��q!��+M�F��V+�r�W�bbH�tl�~lAd�3�=G]�o*��Ԏz��*_N{$)��[�{G{5���H�&D ���L�;F~���tp���ʝ�"��@S���a
���VN�(\v�:����g�0���u�fB-H�pQ�Nݾ�X�u�_uT�L��_�t��S9�_>y�w���e��>�s@)TP�����C��Ap�@d_�'����ΘL�.�Z�1��~B�������w��.�#6t-�d�)��|�:#T4�2W���5���x�q�c��L� �����F��1i�Җi�P��M���J�x���#��_��OCB3����/[R����A��s~�;�:SWK1�l������S^Ļb�G�:M��#�4k�Ñ.�������C���QMv�U�n��~��$Ht�����#2��հ�6#R��D��'pgN�0Mk��*�SJ�dש�˻?0q�1=���� 8B`��n��f�A�Fe5 M�zla��@�c-�lը���]��u�����gVe4Eܬ�m4�>�����aG(�@�ȼ,}Xj�V�;�'�����^��u�,���T̚3�%�"c��)���	�{|07yw��p�)���~������d���"_@E�r��6&����ts_�}s�pc�9��%sT�k���j�/��+�s|�W���#(ar+Y�*e&jpO��2U�+�Q�/љ��+Q�(�~�\�X}f�%�b���B��̢��	�iw�t���4��2�{��z`���qaD��(�kM 3��kGhR^1� k�Z��V�!�nEv^�ϲ|�;R�]À0�~���A��-\���A����;0�	C�EͶ�/�G��#��6�#�g<ǋ��S9@��>���Ž詇�^G0�|�_R*<'�f����ag d���s��eK�X\A%�r������� ��|��φM'��r�����`���
��f�<�7eB�Kk��򞠉���n��ﱀ8��'�z�����S8��1�C�KP3����Y3
,/R)�1�(��Se��X%�YhW���i��IKŇT�~t����c��j�k,x��w�'���:���?��4'�����U��8b���h����-���stor\rPD���} ?��1	��<� �SY�昃��e3t��-�p�z��K�`��C{�.��M��\Ld���g��	y%M�FYj�L��R2�,N(���0QZ=���Z&w-6�F_�a���C��+��b���#Vբ%%�3�x�@�cO��7�$���ǋ�#�4�ξ4>/J�'��������R�mhri��� �1W���~�)nL��[���\��m��KbT��Z{D,(��}r���A��JHovD��'bk�CT<ҳ�~O�.�`�|̂��H����>W���bR�����7�v�7,�4�-����������c���8L���Ep���(ܧ<(��� /��fF���� �L!Q��uڲ1C�e����chN�i�I���(?��Syuc%+:q��~��Mox�#d�,ң���d\��8�Lp�q+li��,/���V�b3!`���_�S$�S�����!��	Ez��=dаާ��'��F���li���h!��AET���i	]U����΄#��@ց�� R�4�C���]��&���`�&-�a���ິ���`~]9ym4��4A��>��t�Hݫ��B��=8B�Arl�����G �|2X:$�0�U�6t�Ш�N#Ę �F`Y? =-chg7���^j�GG���UD�W��-8K����w�Pm�G�ώ�~��I��h<B�v7M�x�ȨQ�\�r���s��4|
@�\i�,�&�La�sP��#.��<t���>�l��V��d�S�n�"[o�M��>���\��Bf��ߨP����@�@��&a� /��b�x�pN.Q�p���o���������[����ln4uj;��4�)�Q�3@99ͷ����8ү�`_�1J�5|Q��v&�5$7��%�,�ƫe� ���}������Ω4뉮z�V48� ��� ��2*{�3Yoʴ�+Fa�Ӑ��H�:/f��r`�� ��X�X~�jC>�Pӭ��'Nw�ˉ	��/qY�{�!@�^j�#ߝf�[�r�ȃ�d��F�Ϋ���w|@3ו*h~`TΏ�>��[�'�E���/G�jui�F��Yޑ�q����	������C-:�V=@�s��wH$^aA�2ҧ��v�������v��쵡���$M��0�arJ��vL�̊ue��LkL���~%`�\��4�mЊx�T}.𼂗�p����}b�(�Z���uEB�㼃Byn�
D��p \H�E *_�Lgy�	��0�*%����LMy�����+F��)g,lWih��2��z��!� {��ADlH�;���:�sCKB�<Q0�l�����$z�MȞ?���&{�/w��S��7�@n*%����(a��9�n��J������O�c�²�&Av�B >�t��i�#p�y>�C�g#�W�<�������P�|K}EW�+�o#�B�Ha.�
�PVe���(����V�B�[�g\o+�C�9�L�<�ý|�_%s�:<��Fca>�<�a��:8%֊��qv�%D�Vo,���7 ������f2�ߗ�����9#��lhf����.Ŵ�cN�p���{�u������b^ ��uvKO�j�YhV��^C�ߔ���tB�9�҂���WDdk0V	�O���j��H�8C�}��{�t�"'x��o���ز�>�\X��jo+Z�Ӷ��hw��ɕ����1 �P������R�=�=M��`�L��OZ���1�MK��>ĽM�/2{	�#�T=�,j^�0��(ژkj�"���ëɰ���PyJ�������u77�>y�Z�3�����1�P?�z�4�[�wk��Ň;�(˂� �!="����+
�y �h����!�����5>���Ps12���׷�I�b�-���}=�N������?�os�;e��7�罝m������Ͳ	}��1����yE�TLE�%�VH*���/"�ո>��*8������C�>I  r]�tj�4���0S�P��M5}�D�Lv���X3�9A�CQ�|��lP����BG�Ѻ�[�yjI���"����ç��nϵ�kd�Cb�r~�Ҿ�#.?�&�,��w�l;ʝ	�\{��N�4n�>�M>����"�Zpd��H`b� �\��N��1.� ��,�Ø8�Ǜ��f?�j��4�O�%����Z�^��npI��EV����;���.�c�zi+М#���nNcр����NU�<��'����JFm���)��T?^�y<|C!�̘4&ÛMv6\:q 
��P\ڥ��r���aO�����}�U��r�v�G𡁈��P`%nh,��������5_7��q����W*4��5�|�{��������P�	L��	�<��	��ֳ�56J��E9k�#�lK�Eb�$���X����{�о�2���6W��p
 2Gs�:=�jXZj���/�Z�*4�^��ă{��c���v-�$��d
�Y�.�����Zf��z��e��V�#�M�)Q�f6�cf���uV�����;�1�w��\����
����$a��S5�ieF��@�ˊ��?���#
b<oQZК�P"Ht�tHc��66~��dxغ��������A��1�:����E%'��ҏ�2h,Rn�TEB�YQ��T>�a��|Y����Op�J�X^��:8v��l�l���;��g�ڌ�|o�*�`�TB�ĺ� �hLu���c�`���lr�?��m?e���r�<Zb�W�=�L�����/-�f�Ѿ�؜|�}-1�)q���3M<�i�[���[!�^Jk�
"�
Ϳ�15���d2npJ�����Lflp[��a�fo�J��!t��߇M�fJڝ0Zo��~PN���̕.�U)<�Ŗ�?�������y �{��Mx'T�~21���)�^vYu�-�Jf�������Ǌ���Vm��m")8^/!��(��""c�������ǹ���M����G������e�l�������x5��w0��������/������:��(F�vlu�r����n���ٱ���#�z1A���	C�_���~}���f��4���]�oHv����I����.���Q�Zsm
/���u2P��Z��s7�ļ�N���9o�&�LW9Pc�5�\ֿ2�����|%,>oX7�U������5LRE��T���	���;!u#�xث�n^ ϫ���±A���1B��
��i�nf�7qVy�^�RDN����N�̧��X�}����p�aY���/]c��cG�K���
�P�HL�o嚷��y��%ө�}@��Xwu�v'�-#ݶ]MW7<�K����7'���I �{���]�5���sW��I�j�p�E��_e�M0�`�D�@�w�+�ѡ�#���>���)r=Q��xr�:�N}��ǚt��<�:L��STH�^V���p�WR��rv��r�)�mÂ�KnNi����#-9:�rx�J��l���ߒB�r��c������q�KG{dH��G�pPtR.ڜ"�����������<��7�����uK��7���:��g�6��Up�U]!�oV��|:����kBL�5����M�ۤ,�?O���F9�J�d5O�R��PDt���Vb�2�������t�o"j1h,���� �c_��I�Uµ��g�Nҳ��!�#�Ĕ|���,<��?_�9nA�R���u�*V���/�5`��>y�W?ܖkC�bFSB��Z�mgcĤ���Ck]���Xz���\��~�kZ�Jq�EA �ɘs3��Q^d;�߻�/��z.���0Wap;3٠5���-�v�=|��ӏ���+�$�^3������Wĉn�ʔ��(Vt_|�'
	s�ҝr$$�_�J�4��K��O�_͋�D�CB��%jE������f��N�\G�c �.�"RZ�pD+knMQ��z���u�����>�9�z�����`��E$��eMv����VO�D�bL%���ܥ4���hb$ws/�Iʬ8�W�od҆/����Fުx�0�,�M��pq�(n�TA�'efx`�L�űp��ql�!ŋ.L���9q��6�s�.�2\~t��ԉ��7�6D���-����ps+����L�!�O:|kZ`1�.b]M�wX��J�R�o��Å�Zo���#�2���<i�;�0��&������F��Oo��\V�� ���rLqM"A��)���#n¥������C�_�Q�� ^�~��z[%��C9P�.C�@�t7�����[O�ՌIp�����+��I�H���/�����Q��Q{�g������]�P!��,hq�0��d�Z`_��j�7ޢf�G蝰���+�q�&�K��y*�&�]����oy�aӨ��^�t����Ĝ��g��S2�������M�)#�MTJ��b��������s���q�a.��C9_)���4�b4��\�V9��m�a��t�t��˚^���+�xV����7k9��D�w��D����m��v/����t|ؠn��wبm��#|����*I�5�,�`Y�;��W��=���w��&|��fC��=Y5�(hݚ�g�A�8�Cޯ���9�f�Bsd�=��}�v:�|��h�D}�h׫�S��C���z�z[�����X%�c�j�8�R'����p�襸1,0�"�-�z�Cm���專s��{/��pj�o�����&}Vs���PHA.qy* t����|��^���׫���_n5����4]�V|V���1�`Z�y�B7K�oF�k�S�!8�ʀ��Ӏ~���{: �0�\8���ć[���>M4>z�N�:�e�u:�sm��&Hi�dG)�]#|����J?Q�j�>I���bfc�`%�V�?G��[��@��=��!A�iWW����������z�%�p���.��� �6A�$�fUԴ�M��mQ��W�t��^rv ���x��
�y*!=�7|�j�Qc�y����\���H�1lQ+JP�l��uX������u���o�Y�(r���g*&��vb�j7�DK���F��*�B'dr{���eڵ3Ph�ݪ��4���E���lL�UJ/X �׳��<n��:����ef&Hѕ� p����;g<��������oӑ4|���df^4��?O�Kl�l�Q�V�-�G����4����[A�,�Ǜ�ry_�e���ɿc�p2oZ��y�������cжq�,���g	�!�J����(N�`@�Zdl���
�PV� ���=ꆌ�@�Wr��e�
̅a��+�(���q�� K�m��\A~�H�蚐��r�hj�+W��mI�^j�p�þr���������x]�\����}`A�HܣP���
d��g@(������+e[�����k��}��9Wb
���� 0��2��\"�[L`5$yN��	�_����ߥ�Qf����ښ��Pf�Y��/��h�!@�2��`�� $3�ª��F�]LL����%ɕ�`��ְ��(�b�������f34��u�D���!��!�<#j�"$9�1[�C��;�>[B�`O��9"��g�/'��r�]N��Пd��8��_�O�	���o �����k\�_���d��&����V�8�v�?�0��!̇ _�Yć��>�+��n⫲�b�v�Ao��v�s�e��ޤq��T�3�K�����Ӧ��J9�O��5�Q�V^�+��ӓ�����go���s�&Re�E��RF�C���k����7C���3����c$�����m�m�:f$E��!hD���~�O�'�����:�X�.#z��F�,4v$�K�My~��(����6>��C{)R`�b����cn�J���1��Ȕ�qx�a�Z��������)�خB��a�L�M��>����B�$Y_yI��m�8!J��[Y��绵���i��ڜ�āK97Zp�H���'��c�e"U�4.���]JۊO"�l�xN5k^�,�ߪ�ҪD��y�|�btfO��|g���'B��H�����M�%1�V�LNO��,U��Ú���{L��WA����S["a��NI�~�oN}9���;�����i�/���{����լ�������, �̆�3�`�����a����l��\���=���,�}�`n!�=y��U!�kE�{!���Ak�r^��X���^��܇�gkz����7B���t�`�E�J*�ޑgz~�ToVʶ�s���1s���d@LrpJ�G�� ޝkp��QWoY1. l/�Zy�X��*@�5/�"�*,��k��)�E��<���lhGupo����>c�Ɋ�k@gh�4�OV���Ҥ}Ⱦ�ė���ʪJ/f�	�����b���v&h��j�1��.��%DDA]��f벺�J0%j["l�<>��r���� 8Ƌ�Қ�P��s���,ǋ��L�ʡ����bY"�b����/�{N<�i�K�>f:ɉ1�|���*7�ˑ\U��N]m��RA�n���M�X�|�֓��N�Nzxpg|��X��;���z�v��Щ$�</`8���w�Bʗ4 8AW|��O��T�T0C��s�	0�ĺ������b���|�.��F8�����KY��O��R��WK�u��nY�=�wВtz"�y�,�� �# Rb�d t؅K��g��l�ߝ�aJ/�@�������컆Ӹڂ�9�;���[�Q�E�@���g������4�E`	��v�<����6?�'�S��jz?�м�%�4�����I�d}�D6s��6OxR�.Xk�hӕ�[;p4XР7�٣؂k��Ú�u���2^�!aV���}^ a������Vb��k	��oC໗!��2EC��߬=d��2�1����i�_S&�Ӫ0�f�	��{��PE�	�ނ���Y�l�3�#��*L��Y/�r�?�˔��まwe"�I�,�#y�
߇ �ܴ7K	���K<�[&b��y�Gs� ��&�g
��Q3�)$�@/�\��iV�3�cȈ������m )�^��q���hs��%�=�ӮO��$���{#R=�1�O�jQ���=���<��`?>����əpKwf-�OF�kҞs4�hn�6���T��/��'�3՜��l�,�>I�?Y�
/I(�ݐ��:�"&��4$xY��GH�dռP��vc��[�l�2�f>��6��œ1�(�>k]6�Q�'
er�2�9_��{���UK�s���W�Q5�=ヮN/��T�먮l6�o.���J�G[���JB�	����z�� �����E����vI2�r��r��ձL��s ��
�1��L�&�;����wB�j��g=��m����k������d�����o��Ws���8���~?��[=	X��r��tPMGA5����/J.QM5q]3Ӹ�nU9�Z&�ڥ��HkK�wT�׫�.��������h�`_Ym�vt�Y�o�
Տ>dэo�eBJKv�~��v?�(���&����TLܯ\ǉ��J��~A�bی�C�oV�H���(��F�o�>�9��-#;b�o��ߓ���#��&mGF�V3x'@/�lXn��:)� ���U�(��FA���,�~��G-��viMVC�ރs��+7*`�z4,�FB�Ί`���%iЎm\ې��zx��C����L�@��<�W�y|M���W��Rz ��э�z�f	���	BQKT,
��@6���?zml�EM#r__�%��Y�-��l���:������}kŝ�l��;�f7.U��H�)-����M��M���cJ��IR���D��9��}�X:Mȁ���V
ج�BF6gK`*�К]���y<�wT��Ew�b�'����D��^-ލte��=�:8ɻ���W�v�������ċ�"!u(��L�V�:lB�w�Й�������nc��FڶA%B�嘀�a�͝f1.y�yl�˵�߀q�[5��9-�)V�����b�V?�m�6���i/A�S^��>� �~!��W�Nh�9c�WaZ��U�o>|N,I�B��>y�]�!�f6��u0=12Vs�N����U����������!�-�������po�s�t#�dJ��D/10V��?@%wi��4ҡ<�ح���)�:�D�H���o�m;Sܑ���C?,�K/��	�2.uMG��=��BY,*+�/8��tuɦ�����
�*v��m���$���՚�"��)���,�qǰ)��$��왟΂��'IYA����"��tS�}=s��h��,�k�cfX��u�e�?��-�\zyR-&�/��\�������`YIk��Yr�d�p
ٙ�s�� L�>��`[��h��e�Y��ư��?p!}�J��3p���U�sa<�u%�o/�|���.<A��]�/Çz��g��<UB�#�St�R7K�yFkG�O
���͛�~���[S�z������x�T�oy<-��z�Vm������/��*��L��w�s��H��|H΅4�Z��dl(Ɉ�X�T���
���R��c�����Û
�D�}����g��^�PM�A[�H�O��b����${#�Ey7m�v��h(�(���'LXn�[m�U���9�7ۄ�rHj�s����m��A�B�w�3�
�ǯ����/�2'*v�ڄ��>)F�F�U�c�$�*㕸�*���t	�6T��.��Ï��֒&f��ς��p;�a��z��Hjab�{(����KbO!oE�*��s��\v��o�� ��o,�l8^g���x�drAiݛ@	9魖^N�,Xa/N������@A;[�]L�	���9w��*V�s�"�w�^�Eߐ�����V~�yϯ{(�w� �a�����씁����Խ[Z��;|4s���on^9Gnqo���\�Ad"�3� 1��W�T[ϭUu%�n^ʃ�+u���Ċ�0HM��!i��bQ��|Ъ���F#z�Uu�
M���"!��/{*m������]�v�=��D�I��=6�\�A'g���c4L�B� V���;���cI.k�g�T�EH�3�V�=�=qv�d�9Xx��	�I@w������cS�v?.�5@J͛`�k�$�WC�d��Ƙ)�N
�����
 ��S)Eή]���i���0
����D|-P�Nq�bA��1���
���s���;�nV3�8��&��J�}� ��*��%�[r;߁hBm��K!+�ë�����'��_/��JוU��Tu���j$�
���i�9ߢ��p�����O�[���+�.��@`,�/�v���~�51�).WY"Ѳ���8�yUűzi(�n��B�b�ǅ�����j�Xv�^i�^it)Í6U�$�P�[;�c��;Ny����~�(�`U��~�cm�N%0���m�Љ�t�>�{�,���W�U���nu��̬�H��f-W>�l챐�x~	�����2Ó��.?�6.����xS'�?K������`5��M,�X6��0�5�����I70�.8��t1�r�N���,��fx!�F4h�{}�Э�{b���^AA�����i"��45�����������j����ٴJR|P�X�.��}6�MY��``�K��XM����K�.�&?�G�(�r����j�r{�/r�أ��e]������f���52���A"�N|��e��nY���A5�&�����������zn>͇�`Y��`^��g�� Hv�~�{;J�<��LT�<��� �R#$�E�7ݣ�ݎ�-GGɢfJ:�V�'��>b����rv߄�Ь�芨�-�w}VX�Fߞ/����>>�c4��	�����p�1Uحϯ���P"��:.�*:����@�4�ʸ��!d|���L������m��:Pw�D�6%��K�y�@�U�gc�����d٫�p�)L��� AFg�*��̊Z��DPK�̘z,PgD�=��Rc��ϗz}��*�ӡ�F|�oG���ӻ�q��_�s��������HB��i��E^������n�	���%�@CQ��訣3?��+��y��N޺��)�8�v�"����2X��G+�Baj������Ho�	F�՚����$���h�+��?r��@�����k�o;��V���քsn�;��9���)��)9e���6�џ��IG���:�ffxv�K�P��&A�����FJ>���s��<��oQ�r��A�?#>�䫩���$�
�e�9�^�~(��U.]��!s���-�O��Xk'�y�V��~��W2]b�bp����L��jj���^QW��Ba/�f�P-n'�eD����Ar<� K�ͥ<V��	M�-�%��*��eȀT�"5��������$f����I�k���rM:�k-|��J�]�e��IR���pj{wȞ��=4�;�.ί<��>�[��2F�~7>�9�+O�+g/,bl�Ug'HH��.��0�^���b��ρJL�؋` ���Ip�mн��
�Mu^d�V;.�&_�`�H���SX�z�jh����F@,>�>�UU��r�� �³Rq������!�Vco�O�z:�_�W�����ەhң��U&�6Qi^� �=Hi@�"��"���|ݴŴLz�>t����Kc�p�!��*�3N���d'�����-ԙ�D�H}4�bSc�W ��yd�p�ϿFH1���n����}P_J�c����*09[�eo�;���qd�РKy؜(~Z��o���4���5�߰.�'~,2\�Rf��c%� �8Uϥ�x\�z�mm��*n�ԧQ�,�u��E��_�ψ�k+�6(d�|�oHO�ӛ��jY�snNA���K�A�2�l[!ڿH�Iq�/r~�n �B|䉳��n:��{�һ�{�7F�i�����rd	��61�r� p�#hR���f���/��#�-L
���Wo�P�%��95��BqV@]��X��G�B& ���R���#^霢�p^�-��j��1��k�oU/����({��H�fA?�m�}������c��[�&Q����5���ڿd'�<�|���~��ݡ�I�w�L�13����zS��F��6���+J�~�`��,�-�t�ID�Y�՘�����9�JD�)����1� ��k0�$a���D�ԼQ�2T*6k|:�N-"��b+�'\�d1�t���Ʃ�!�-��̷�}(N��K��ډ��l6fu�-$\�6��zBz;�}b5WjF�l�M\�����`]B0.����mE��~S̎�4�N���A�O�P2FIFy���3� y��|�,d~��S@Xg�>�.b�͘�
.�������W���S�nr(p���u��;�\#�,F������ې����2��s��$lg�z�'��A�ŊbK�ȊX5�炣9�T1�7�N1���I��*銪�qfQ #���a�oUְ'b�g�4��[Y�?�g(f��g,CC�@l�O��^��d
�WÁٹU���w�>���s�QzD��m�wӺG����F�E�*��s�V�fѡ���,��M9|~�&q��!�����x�i"�8l$��=��T�Q�SN"���f�]�
?���J�X��ap�?��n����v����@[,(�(����¦���h粑���j�J�y���)@�D�Mi��/�v�z�$O��.�A`���Ɯ�"b�#*��J��I��:��k��-��b���Ϩ�������'[�+���p��g���m#�6��Q/��t�uT�qO/�����k��'m�=9�����>�\�	m'(��0;��C��7�bla&/��h'#ߠ��!o��	�7�/CT�K*N6d�A�=nHn*q�J�ԫ����S"�K��6���^�������qہl�H|�+;��1���)��3��cw @��Q�̏���.�EÙ,�B���@E��[�d6���]�����.�I�.�(�~Q>���z���ˉ,����h�@�5hv����P��T�&Hɤ�3����۬mm7M���#8Cr:G�:'�;�3j��N���0�u�v���
�g5��ב�nd�+X,��<Ưk�(yF-�.��C3%�tl�$p���u�)�I�]=#;<��7G(3�K��C�C�X�XܮI�P��ZN�;l�~0����7M��Bz�zkc@��%Ը�b�r��g�[��\ �5J�P$s�{�����ݳ����(�2	�I@�M��7�7􏆜����:�߀J�4I��eP	�T�y�_�)n��Q�ߠ���B���9��-^�n*^(�.R��Sm�E������.�I"��[�+�͘�qwN}�{Ҭ6�9?y�"� ~��5��0`��g�3·3B�T"��*���E�E����<�VB� ��U�[��y�Y[\ҽνD��("7�_7L!��=+�[�3n��c�4j����r��\��o�jnX݅>�x��Q�z6*�~�QO�ƥ�����iJN":�K?�[V��E�P52���j=��ʮ���ӏ�b�`}�[-*1�˛�%r�8ி�f�( ڄ�u�?/�Dƪ�3f�%��)���Ex'��+��������?��M���y��Σw���{f�+��QQ�����[���6�SD� ��*X~`�#ꕺ.+�*᪽�!����לIa���C'gK�>���N�j�w` ��u�(8��v��`��hf�G��xf����C�<9$&�U�V\�1�����9Pv��^�M��^��[-�n�)�ן�t���������Z
�aq�f��Z]>�?_���_��|��$ܝ�g7bÖ5�/m&*̦c���s#�f �/Ѩ,���'IQ?,i��Ƞi��v���ޘ�ʆ�?0 $3�/UߦP�d���7�ŔF�rr��,M���"�S]��qǢ��q���V���`6����BS�/�-x���Z��N�)�L�f&`�e�P$?�.%Q:+�ȣ�
#����J��^�h�����AO|<g�;�Դ��vXh��j��k��kC��Կ��cAl1��9�C F����V:��t�����vr�a��B�4/��D �"�+��O$�t!_��p�*]� l"�SK��ދ�O�YJ��n�WaQ���PO}����P�h��Ʋ�6���-JI���_H�;�9�EM�̻uQ���\��M�Y�k��Rɕ���<]��?�@�_H�QO�	/��6����{]ȸØ�q1�|�W��F��!F�/���|v�~�٫�<��KO����{`���E��Da�����j�2���,է;<��p\ (�S�K���i������1Á"�ɨ�҆��dq���R��}0�@@N§9ɤ�Y6��,��	-� F��0G�t�7���%�A����*��L��1�z����֚��]xa-�0���okq��^HCa���/�r��H�k��4"/s4挒�.Ѷ��F�\��"�B�K%/<'���nH0���@����:�L.G�9w���z�����g���%��Цq7kR���{*��Ff��'��"VB4�Y�����W��4��h�w�S��y4'V����;
 �4d����%N��a�Ƽ^�]��ީ@�] � �����% FZ���^��?�
��m0�uU��5�ǧ����<C������O� ��wvࢩ��E�`4*���5�A�~�|�_ȵ0�E�QXz�{�%)&V��-�)!Ƌ�����a}3��[^�X�$Wg�rM�G)�|9�;�RN��,"�U!N A��S,{�<A�wMП��������`�p�T���)$�����i�e��e#\�S�K`�=�v�T�F(���#�J���hBqB/FT�U`�K�d��1����" B����rbJ
!cZM��[C�*!A�e���h~����c�p|��c6p#`#��?�펣`�s0Qi��G|2Ps)<'v���g	�&S(�&��0.?'%���J3Z��H��U���݋�%5lk�X=�$��G�4��QE�*�)MFe�<?��=H٬��*��a4����1Zv�I/~w�����bd{��6s��`
a��)����t�4TǄe��,�u6!���ma�N)%r M�Kwt��m�����RP�����S;���{ν����q��'�[	�6��Nx �򄷤l�F���^�����Ɩl&
"d+�/<��|�7�V����Ǹ_��F��eV��V�Uc�&������������uL�r�|��	d�J�B����H����{��ó��4�6VF,�(��6c�w�M�6��XKh;`��o�ŃtZIK���B>1/_��|@���)(s�rR�����gZ��	I��;���g�|�sX���Ь��"" ���0T۬�(V���k�rQg�F�,+ȒȢ^i�=��h�^C��ïm��d��;EӦ���]�����R�0��2�Ʋ{���NǗ$���rs4�BΟ��-;�2�{d?�t��x�5��.��(6T��� �� ��R�Z��S�u{-SN%+GRX(�l���EGp�8�u�D��>�|��"1.��G��'������� '�p�9�wF=�;;k�Y���>��$eW=<�#ӁJJ ���=�J�eǥ`�t�(�Hj�T��; �ӎ�.)9�7�~���*�i	�.�m��j�*�&�6M�s[b���w�FJ5M���-�j��%�Ys�}K���=w��ƀ�K$�:0��I��2ŧ*��8��=Q���!�gx���m��%I?�U4"+0V��j@�b�ᵐ��?F�(���o�-�ay�{���y���q���I6a��@ק���SO�o��@Ig}g�D��V��ۆ�$.;�;��B׎�?.�%�� ���_ˡ�L��L�g�q'-1]m��[q���!E*�%P� ��|
!O�pf�۫��p���Y�.$�g����HZ]
�g�`�=H"9���2+
�,�y	ڝ�إ�S��]9������=��&�z��֚����īܺ]�+�ř3��IX�5�H[%A�(3�f������2fޫ�-T�k���t�qo�t����,�P�n&��q�y���#\	����7�f\9l��0���&�Ɵ��;�|&�^,�c��(Ưd�`���h�C\�K��o����iPSq��h���%'�S�Ĵ�Ӻ��c�c"6���팚�*�џ�U�B{M��GcR����e�.������ �_	,��W@`\�e#�ض�{5������$j�#ɤL��\��~�({��h����PE�3��tP�\���Ms�')��ww�9�y}i6�'Bj`
U���eb��+��-�&�O�_.�ϊ��w���bY:�Ş
$�3|�Qy';ް�N]����Ks�w��Z,][�0�Z�T^�B�
���Eɔx�w�� X�|M�U9��L���X��
�I�*�Z�:��}#uù�Ad�������4�n�P{�!���&�Y~�sɠ`sv]SD&M�&�s��׸�	 �vg�Ze��oP)
b6D=�9d�0�O]�O�˷������A$�@ݒ򠬐�a��)BD%��ٺ���*'�Ks�P[��]�M���FZ��*����n15�A�kd5\��r�$Rb��ڱ�8�,�{T��WM)���U,u���Kf���"9��\�1>o�a��w���H�G����w8;�8ǏݔK;[��#	_.X|������@���!���1sD�[E��|n{�b�;��������e�۫q��-��V�!�$_w	��<50FW��${��]�U�em��� ��W����N-��z��!�sY�܁�w��G�_
ޙ,�x5e������zҹ�o�TS<����]BR8��!��zu4�q%��bL�hs�#�]8����n��Ou�@�]�:T���Yu��A�0B�(X|���S�#�Ā�.}��SY���1#�~ME����Q� �G�pZP�({?'ʉ���G���,.�!��h�X����?)[������'u^�l�e��M�c�+���>���6�%����3�����K%(�	ܹF�Z�qF/��q��mo#�3�Ĝ�7���c"W2�؀�$����%����CE	͹1ns�UG����<�=>�w��c�.�?J�;�l�Ƃ���̷@�o�	��s���&];��Aæ9Ylgj3F�k�;�*��gǥUs��Pb�?.��"f���m��]h��k5���<A��B]��w�f\#�)�b+!-��k$�/�Q��Z0���%�4Z�Fs�ZD@8�ɲ���"�!����%Z�����+�i�qÛ��L\f����I-0�.`v�c�r����܋��xw�]�_���ʯ
K����W���"=,�rd�����F��q���9��l@��i�����\��9f\ދ�K�~C�$똈K�.�~�!���6Ͷ�t-r�6��u�s� 2S�4k$.>R�(�?�x�|Ht��L#�������F��,�z+!۩�R.��)�a�-Q�g��MF��.��0�n"P2��\�T.M�t��>��%�"�%P��1JG3)��>�Uhi	�gP֌��*U%WƓ�.p̚��)��[w����]���6AVO͇�ԫF��K;>Ӫ�_HP鰢if>����#!p�����EҼ���{�;���T?o�����&�#~�?����^�U���3Ŧw���=167�K&>,��.���asu��)%06�`�
�����:+���Uڃ�W�j�6��5$�V2@�n��JI!�jn���#w'b�0���a޿ݏO �,(���!I*d��Z�5��,m�FkA�����6�ْ��mx��.]ӧN�4�����$[�ew�GR>h�E���GC.qg�����cY�`N6Ð��N@�"
�>��@ ��/17_a����WtK��>�Ղ$�YƂn���z�Dcc�T)v�9]n�{�1��Xtf	¡)����'.BS�rҲ\s'�/q�=<$�(�P{O�B�
E���kROƏ#'b�o� +�F@:D�Ԟ^;X.hM���� r؈!6נW��ߖ�@��=��qe9	P\$����^�U��s��N�AO�%"�]�<��T{A-���Kv�	륊H;�ξ�ϸ/|ʍ<5N�c`�����,&!>�B�E��x��Yk �ʨ�C=Z���A������s(&� !�My2�)��sQ>�V)t�d]��	�?	:�@X��vi��gڐ�y�C,�p�o�Q���R���E����,!�	[-�7�A��P?�e�S����T��P�-oLf��#�¸ڡ�[Tȼ��d7_��6����Xt���3IHN�S颤2�/�����
?��/�����m�7���b �����������RO�	(�|�.{�01�^`<3Q}.3����`��ı�#5�tY�K���,*�q�#��؁�}?2�����wH��Y �?W�w��%О=.g.�z��+��`$��A�������1�t�K4i��/�ȑ���8�lw��#��m�_���v�c�q4n: �%T+x����A;��Ϫ�K�v���~�
���R���Ƀ��B�`P��k�n8��N�d��)�Ir���{3�I�P���n3�w,���$eG��?!�:riX�v!�����zQ����er���3ꅜc����\�
%H�~���H�~��C�֓{�u��E�J�}�����1�l�`�sԩ�FJM`4�
���x)���Sb|��Ⱦ�[c]�O������;5�h�a�b����UTw_i��1�4�����Q�a������9�L��xvHH©�	�b����'�������K�8��3�'�,@�M@(},u�;r�p��cg�p���K�x��r�r�>D<��o�|%����qn�������@��^- �+Z��^��_ב��
�֤b�sl��XA���soZ!��,V�7���M�W�e�s����bG	�n�L�s�no��tz4�ڹg7��O5� �3z9�/j�7e����F�~�6���S�j�-���xo�vl]��-��R	���p�Ô�@����j��uk�hQS����i�)�]��\K�s�/����C�~"�*5*�)E��'~Q�$���Z:Et���p7�p��N�J�U��p$72&XB� `�Bk�"�`~��~tFx�d� D��9�qzu*�T�a�E�Ֆ���?C�E��� ��\.����aLd.���0s���̠ZyrJ�uJ���L���,~�N���1Y]�w�5��s�I�,��8 D�,��:WG�1�S#.a���Գ@����W��z�Aո��G��Ɍ�N;��+�?�.���.*G�3(�l�, ���rXo�y�"ゥɼ�"X�R� @��uI��E�Pt�����RZN�/ƦI"�\~�^����ë��Z��) Z�; c���c�(t "a!�`dx��XG`F��O�|�EW�'M,�M�nU.ߠ����U��
�IUhY�A�iw���Iz=���Ɛ�Ȼ�ֽtG#A�IS_�+ۘ+��0�H��?���J��o����}�S\��m�(�u������8���:��fZⷐ&>�"����7oMd���?ZEj
B�j4�}�ݺ�5�	��]���AgYL9�4�X�A�hHh) S�;K�F�$�G1��5����ڟ
8F����l$&>��Xr��@���#ڕL�����z�s5�v ���s�|�m$a���$��Oҝ�7���,N��:�s'�
�+�
�g���z�r���S�F��g{��{�n�oM��>�c�$�@��g��a	L
W�-�=��9ҘF�(:��A�;W�\a�ϐ����;��H����?����5������.�3��p�H��:��uI��π���}I��'�)!���t�_���z�
�_td��6<���c�=@'�:�\��̧� ���伞�G��k���d���yR���+F�������P
w��E�p��MzGˣ�˰������)���՛���Y�:X� �%PF�Pw�����U-���3�&�0.��oK�NSM^<�r���I����uz�7W�.��:����;(	e�\�V��T�g��n+M��k���Kc�f�Y�8�c����}�iŇ����,l¡����㈗��C~�+�L���S��5o:�|\�t�M7����!�J�r��fO�GL��Q��Q�M\��Ş�8�Q��B��:ƍ5'aJ�x@rm���Br���(Ӈ�y���Y:�g�Ѯ�'(�^��0�u$��m嫶���0��!�+4��D>%QLX֒�}S�^L�_��|5��-�ț]V����۵��j{7^$̙�c���8w;�?���A��\�H+�՝�%�n^��V#��Yd4�ܲ�"[�f�	������:��#���F��PV_�P<���O=��h،*;��^��:����b�w�A���?�=lhp��ͭ�����J��f8o@*�⢍���#̂܁wsj�����D<���W����ϫn�B��\�_��cQjs���z��C ���a �|x�*����'��CF�Տ��u���>�e�u�G�r���U���������Y#��ن��Ҝ�yz|��ғ��z���ܚY~���Q���TՎ����`�l�,ظv��
W1�F'�����M(Ǜ9�8Ck�Q;�Sf�3p�qq
!R��N�U�`���4�E5=:��C�&f��62^�~J�u	��p�h�m51�6Bё�p"��(F:!9���	�5�YE0^B��D���!r�U�`M����赒�{8�����Ht�����
�<�z�?�߇֬_C�+� iĔ+-\.ѦO�[���rah6j6s�E� ��Nl�4D��v��u�A���u���-�O���f���̆�H����D?���\�-��A�!T��0c�j/XZ.
b�a-7E�?�E�v�+�+�8�l(�x
u�Z6߻h����8(��8E�1�[0�Un[�`5W�;+�"9��#׊��q��9��,�O��z�]<a���ծf%��h�9��N�Y*�e?�y�kE��{�O@�}'+�j�4������
��8�>���qE����?����$�7�b���~cާ�C�3ҧZ�l�_��v`�de@� �M�TW�ˆ̨b�Ke�eM��蚂#�&!�����KF_���]��5e�|�8��:	lõ�r�Ι���]H�-�7���!��e�R��
T�,�E@��ٝ�˚ϲ��y�ͅ!:�[7f��}��x� ( �6���Oc����Ob�S��>S?[�������
�Q!��V�q:qId-���2��b�5��%8�����pG�*y�d�P��P�Y0B��q����Б��e��V�R��&� Z8�9I�����%��֎o�F���ʈ��-�0s?����ظ�t}��P �J3����fbf�c &�-�@��G�m��'���=yPgW3*�Q�}}�F�v�O�f��Y��ib�-A��@��DR)~2)�(V�K�8Έ#��	D؊��	�I:�l���M�1��o	��l��<�*D���֔�>v���Z��p�SI�ި#)>��(�¢�U�C!δ������&�n��4E5�9v_d�:��K9=H`JC	���bO�}�5��QNO���M,��H/�����gޮ���]��QX�Z�<�{��|�µ7�
C�E���vGE�^o�L8�&z��+�j	,��$�s��*��V�(#��(h����z"e��d�9�6e���;�F���[/Xl��/*��r2-���\�uD�٦w\�_�����&�D��,	�ht��,ו�C�)`�����6B,���O1�5�+t�<�>�����=�l����
i��Z%Pl�?����&�RyE�m&��8ցtGz/�FwX*!������v�V.�_>0͙�P�'�8��(	���?mө ;��S�:ﵴ�g�bg%o��_`0e�WIt��`R��p���<Tp���W,P�x��i����!U1��h��ٝ��H��r$#��G��.(�`��t�(.��#{q\�"�цQ��8b���������m��:���.a��$�)0��Ӯ1��Q;?T�)�!\��� �>@��&���<!cV
�v��\5����E���m��I.������bj5o�ī� ��Q�{9�a���7��"1G�{��xyn�e� rw�L����1=����f�ZE�o�[�,"���a��b(�:��;�A�M��hb���r�*�̚�'�y�ސ���ջ�x=m#��U[�Q!�����5yutD[�:>ŀ�Um�d7��n��d~W�TOr��Ե���M�"����*��K(�T��>l'W�k��R�I�l�1�����j.����.ܢ^ȵ�@8���W��(�"ִ�����d�AsYBd"I�̻f���,�R���	Fd���t0�Y��h^͇�2`�Zmm�	f�*� F��nU�ӧ���OI�<���7�;Q��)��Y�0���iT��OM88*;�T�Y��oE���?w��������%VЪ U�G������ qr��s��W"��NB ��o�J�^i��Aby\�"QWPI���O���ا$W۽�ݡ��5�w� O� �B^an��c����>�+Bc�[�7������*���������\�4VNK����Ʌ��e�Hi��J�f���=�V����`W�F�dï��s�)��N�ʋ���p��}?�Q<V�5�j?�%����J�7��8��s�y72�d����
�/��Y����Tn������*������6��$U��6w���r_@	�{F�\��#����X�R��|�+lT�!R��JvO��X��Eɟ�폤c�2nW�����͘f!F�ε���9!S?A��=�3������uC�-����4@wRSŌ�x�N9N�o����^�ѳ�_|F�r|��p�\⬴N��c��22�-y���C��Gȟ������@����S⌍� �eg�ƺu��.,0�$r}K)F��n�:]�HG��&+����M�=��*��	;�'o>���-)=��M�2�����X�܊�S�O��� �-��p&��r;*��'!����s
PU�b�0Y��H0�K�+ޛNX���U;�[��q�>�5�.��d������c�W'��@A�j�
�q����3��������~�M�a+�lv\,��RQ�3�˹J�L��&D�.������L�Oj��x���M���z�`rS�}#l�+*md���;QST�v�_R��Ҿ�ڸ�U~�04B�kl�oKW��[�j�>����'��^zw�/��p^"T 0�|+,� D�=*���8��#�z|�P3���|��_��9�z�q�x��������h��D��`��� ���7槻3�,7U��U��*8ݴm��s�)�����i�> �����t[�z*`r��B���|��յ"0	����W�^VK��"�vU7H�R<e�B�`��k]�����߶��۟P��L�Y��c~�R��)Q.d�*l�B|X���Sr+�^�G,e�
ȏ
�3t�{{���[�|`!(cǡ՚'�(�<�̪�K�BL/2+��������ԯ��C�35�(ܟ��B��؛19�\G����=��y���m?��N,sמ���ϛPL�`0���s:>N����C���9n4~q�P���R�%�A?h8���uձ��W/����y.Ezޘ?ۗʿ��r!��k��L��!�Ij�&Ж�s7�?��ީuB�xD|us����n\{AGj��V��w*�&���X1�Hh0c �<�P�ƶ>��	{˯����ί�����@�ҧ���>�q�.:M�I�2�*(e%/��˅PK����^dϛ�+M�ȵR�����&~�!��'�f/I�k���/ u�,(=9c�JJ��doA��3�o���� �7�VnĂJ����W塦Z �^���G ��W�~�Uޠ�	��B����ǟ]���,@^��@�LΈ ��"Ma�+���C��A�MH]o����;< }}�߬Օ�<�N���Ғ�Jg�����&��}�N���u��ϙf�t|ǁYp')39^]9l'b*��;�K�'�w��C+��z�%
B����D<0�W驋�>��i�#�Sz�]�y+ +Mn^���2��H>���)g��e���$Ŭ�ת�U�'��N��k����#WcN�At�Mw�9B�Ep;0H8ĥs���_��SB�d�"��<*�ԓ1b�����e�@��V�	վ.~�0=�RHW3�܂�6�{�������U�H�9�3w��y�޾̥d�f�%YHµv�B�JW��t�҆ӣ�c�\��brZs�0o�����I��G�����ep��I�e���4T�� �p��
��� �.��ȡ5�HO�*�d�B�>>Y�)�Q6d7K��j#��N/��`l��>�G��c�0a#~�(�J%�.�l��U�����ԡ���!�۰xx��`��Z��;=���7�����f���qx��I�J$�P������5+N��
�"2���+����,A}�F����*�14��@�����sJ2�=�#�a�@�nugЭ���[2���n�
�?�}dar�4}��of|�Ry��w����YY����p�Ս΢�82�_91BXN�uU���ƅ�MGokY3�a�'�;��o�)yAV��b�':�p����S ��ry�gT���U�$/�}�7 ��jd=Fd��m���y�E�m�5����%�*8e��a��G^��� gxzK�s|u|�h��'R�*���-	�`��#��r�{,�F����؏��1�a���*���i�(���-��x���W���Ǒ���+CS�����?85`܍:j����ak�� S���v/�Azy��e��[5���f947��9�0�˒)	���I��  À��j
�������t�����!�ݭ
�{��k��h/\w	�ɲK1�9��=[��m��� �,�`�]d�=o@g�zg�i��M4�aO0J�����	��r�2���Y�E�A
\��]}�JY�:Qh���霧x�1�TH���)M�⭠��}�~�:j�9�f��1������Vh[�Nے=����`s+��X|:�^9�܏��g��
L��c����"R<!e�z�s��(H4X|�'��@��t�4V�2��|5ܳ��[�Z�1��mA� ��(����o�,Hr���,*����7�w�B詤|�F4t U0w-��3��Z�[�g��Gv��IR�wSC_�i�ޣ/1Q�F��-cc��h�[q��j���5���@%��#���L?b>�²�n�˒��B�¾���m�A0��0s?�%�W-5N�0��t	d����F�����G�/�5�bv�c�*"�7����.'�ȴk�b�X%qÒ�dm<$颃2�����:۱�q��7>�!�IQrP�RuȜ��3��r�Ջ')�hB����aA��m�h�,��+�)���$w^lZ��r) �v�"m�nV�����]��_a��8�U<�xphi?�+����K*�ݐp�/X���lH�w9aq�A.4��Q��Θ(��NX����Z�����QQB��:	���6�'jF��|H�܎��rC���C�Pg6�A��:��� /�f+��l'4�R�='.tF�g�1�Q��|��gm�3mE� 3�3�Ng�����⏬%�}��?!���*�enl-J%���9m�š�b���U��>g;�]T��p[�X(�>˳�b��La@���z�L�E�)O֛�q���u)�K�BV���<?·��2ى�;�$��4��t&4�����z"
;�kKԠ1���?w����=Ѣ��Ḥ����������6�x w�\�R�p�BoU��=4Z�7��������v){��4���"��SJ��t񑵀)�U��%�����-��aȂ� #�K ���^�\MN�~~Q�NJ�]���r�����,Y�K]���-�X��Gc=`2�7�a�	������1YK�Y{kj3&HH��/&�6�0E�5a, S�1�7����2yg�d�O����O�F���]��ǂ3��S��ţ�]��4"Ap�[����>�M��$�2�V�g@��>�,y�����p&y�X�@�;�����Ę`,����#!Ax�vp��d��d{�Xi�G�^srQlz�̌J��Yq��Uq-����\F�n�l$���s�4�Q�x��h����W�i}�vf��"߇���%�����2g�/�<�Ә�PPR*a�V�s��Hd^pW󃗭j��v��[<�:ᬒ�'_l/Mղ��'�G^�8�R?x��d�t,0k�Mi �iܱ�����F�s��j0	���>��xVϻ\?�%/��fJ����{z���C�%�NKBZ�a~M�ip��)�����D�O3E�z��I����^�Ù�3�<�/&�:f�9��|�o&�1�[�ENs.�I���׏v{���sQ��ɠ5[�M�-�M>k8b��C�3�Xmt1�����U���u��,���R|XD���N��O��~�6~�'Tˋ�¬#P��L��P��(�9f�c�v}JL����i�	s�;�"�Ps|N���8IT:Y��SX�zr��PL��a}z��-@���٦�[KL��8�^S�T�o���e��YT���;�?�F�-c���B��c��`�2ÉO�$r�Ӱ���23 �[L.�8�6 @_�Drܦ$c��v���љ�h�n+:�cv��ܞ��6�?�_�H#��k����r�A@�J�$��@Lj;�zhb��G&���!-�O@%Yf:"k=��d]+��6p|�ޖRρ+�ӡo����'vAAo'�;Z.�(���E�!�������t~i��F" y4D���q��	\���4�Z
�CZ	�4,�W-D�ȱ�ke��-p�O:$I39I�F�����%\5ĕX�}�E!�/���,!���h⛌�������8��?��i�<S<#�4{��CaZ��A<dܡ���J�b�L����!cp�Upi��YQf���DG~Ak��6��i�+�ۋ��ȉt�����6`cg��S�8]ν�Z�������<���<H�8�y�>��L��:�5�tT4[у���?��lh��NL0`��3������
̦��4輧R4�ӗ��)�43t��$�W��i4��#����tt�zO1��L�k&C�A��x��P�sH3��P��E�.��]X<.$�OA�F���?��IϹ��ō	U�L'���
^ �J��sn�ֶI�W�����.�v��ڵ�D�ȁ�����P]@�n��oEI��'u�<�	��6��������	ʰY���!y(V�}�_�9$��A��1в���~�=��^��r�rZnܪ���2��H�M�3OXÕ?���c��M����J�Z9g�H��Q8��q<Z�����p���M�'�J�܂�pK�E��N>�Zc){�!C��\�6�ph���)�xx�@WݯU;<�w�<�&9�{�t9J�86�	����/�j/��F��~;��`{��:N��rR��b�#tI����<��P�E�e���7ȕu����%ӎ�G�Dư����PNi����N�4"u���yev�%�	Ź�W63�M:�����ɟ�@4�)M�ؚ��e_��1�f���m�09�mW;b��(a��Tm�x+�X��Y�CQ#����0f�/t���E�y�x��gX-�X+�!2����QSx�p_��Y,�� 	W�D���K͑0��;�i"�#�@�OCyp��F�RN{G�bQ��#Y�]�=XWu��qK$��*&�T�c]{�yx�	r)L�d�9���:1�	�g[8�^��y���QdaG�h��G�~��CBGۨ�Fw*��(;�S�%
�_M�]D�s-_��l��NN�vw�[�$F�h#�{���;>�o8ǷH:���'|��ЙJ��k�G�y�E��M�c	bQLգ:߫ҙ��r��3����������;W>��殳GJ�`�C͠@�e3��J��!>u��Ԃ'�]�#�pt�:�}��u�~�RX����7W���J��m���\�x[�cxEK��sB���4��
%����ᘟ�f��*�V��G�5���w�y��q;������Gπ��CB��O��S@��=Q>^�d��Un褤L!�B� K$�-�a1E� O�
#X�l�(������t�z;J����B�0�YG�r�uG��6�I��?���2s�og��@�&C"{��{f�-���`)ר�z��������i���)��(t��@b���n�������ٓ$/qQ'w��S~�X�%i�e3QU�Lu���v�T|�<���{~�<".�Ar������m�ޚz�[��	8(k �����4L���[UcH�z
�g�#�4b���Y����R��Ds8��O�ǳ�@���8������T��J�e��d�r(����X�]+i�+<�?D��ZߍmdK�o���u�|}7���n�=Բjs�^�E��� twV'�ֹH�ԴJj�
.��8.K���4���u��.4^����{�F��t�ꗝU�s *[ؿ��2^q!
��Ln?!z�6�(�iAD��P%�fIw]����mC��>����e=�F2u��>�*5����M=5�3Z��|fţ�D����|ʭ���b.��`+8����A�NN\؆�w��U���!�e�F�d�DJ.�$�3��M��g@�d?��4�Qp��;C0���_�����_Ф�4�>�L��F�d���#O�[}�
���?:8�zN �d��K�<V��%��C�|��d%�U�݋��������ιŲ�(�J��C�e[N(��G�X�
|�Y���Hn������q������ÚW#p�2_d3�6�.jX\���cs�w�KP����q��1)>��J�a����O́��Q���/�P�1����}*��eY�u
E�*��}"o���tMbB�a	}�Q�ytSc^\�~oY��F6�X�!P��|)8Ha���7!�!w7��<��Zg$ItՉ��v�Q�ܾWZ��
V�B+b�� /,�����V^W#�gUmJ.��)��Y�-����q6�c0Ҷ-���n���m��Au�����M5�����������Xw�,4����J�p�D�W��'ʕlm�<�ߵ��p��}=8�@�$�a��W�X�J}�����Bm�"���k�Ծ1S�'è�x)�����*�s`X29!U�eCVqb�@L�v�ㇿ&3N�j��`���g&Ck2e��|�a��,=�����.�z����k�Ldt���jW�(��Op���"��+���ף�~B�rƤ��j�l:L��;kL�f,�aOj�i��`�2� VZ���]����h��(�z�X����+5B���db5U} ���}�pͲ����Yi�?���ˁ�m�V @��ʌ���3���
7t�����V�s����.�ϲ�w�����Bq���w&>>&�[6Y�w)��w��l4H�`)97G,I�Ӄq��k�K^��'a��̖u�U��64d&n��C<[��4�WCS�I�jur��؎"S^�q�a�*G��$o�s���{�o�`�؟��ג@�6f\nG|1c�|��=�(�����g��_q�"������^�!5�=W�ͩS���l�u�����F���.��ԻN��TQ>�:�����ơt3��>�`�r^}�q,4��S8�g]��N��]eU�Ӓf�^Bs�D�#���Su���irQ�?3�5����]�HŒ#��BH�_�/��/�[�n<	��T���QCO�%���WpC�k�H���^~��	��4�)�io��:�q�*3Bb&�Jd.@�L�� �HI�6�~ym��n1A���z|�\#�Dr�S?�'�M��|�ק�y�O/��N`ˁ�h��c�-+h�·�d�
)�����Ǆ{{"���;ub���D毇��JGY��C�<��ЧA.��o�� ��{�]c�Ψ�X��܍�RH��ң���ȋ��5x�w��?�L���Q��a�&@�qU�I�����,8�轨?5.�j�b���e��1o�Tv=�[�B�X��p�J��b���R�H9������bE�L/)��m�;���X%g���P�:�,��u��KXᮁ\4���FD���~:gP�|nk��op��5����p���%%�OZȔ��a�#�L�k�hG��0�t��J��O"7�{5��б)B�UC,�teq[�: �Z�.��@e<���AHE�J���^r̐�C/�!��p\)o0R�ɴ��{�W�cn�\g``d8�5!,v�r�C�.�j��mv�Y�%�Җ���W/#�L����O-ƾjȢ}+o��-���~CD��h���M��\g��Ē���Hl��F�� �)�ݡ@$ �}���q5�};�*�{O���ѽC��d������Z���%�k)"=q2�}�Q�!���.�zm���SK?j}nu{�v�W��Cؼ�i�����+=3��l	�Nl���5�b��.CSQ{Y�r�]	�-c��tF��J����؁p�)v�x/[T|X[��:���?��#��HǙ|��q��j�q~�����@?j@��dP2R����%�Mw�]��O�8 m�X���dЫ��*"G�:n�7kBG7��6id��cm����|����C[w�O<�<�F;��0�{"����ff����sJda�4���fb/�8Y�n~����$%zs?X(���-eC�ذwRm�����vI ��W�ȅI`�����wa�}OA�>$2�WL�GB_r�K�h���Q):��ς�z4�)
�u󖦘����<(y��Me_Y<����a(��^��Ǟ�Z���&@^QQ��D�N�~�)�o�>R���V�ӥ|Yrc���WL~!<�*5.�f�s#�n/[��S�/��n�Z���n ��Z${T��IKe��
�Ѭ�U|9�[��yC�]|	3��;r�B�K��J(>�Y:w�mJP�\w$t�_�y`ٸ����%�.��g^����HD�/����ue!g+���G.�3�mr?��!.�^�+�@2�2�ɿ���Ϡ�a�KM� �Ðm�i}�`��g��J�F&A�^x��!#q���#%W`�S�cP��J;=�C����e�"v{�WSLuR°�4N�=p�ʋ�d?�e�����/��B&�.'�!{x������!�`��(VV:����qN��D[@�qD����l�b]��[��*�mQEB�͠e
-Rʔ���h��9V��f��?��r|��}�
����	B0+ٽ����K���!�-;ƕ䮖%g��˧�����Z?��������zҽ�NX����y|��k��Z&��m���S����v�jQz�i�9��~
?Qg�U��N���Ǘ��=�^x��>;Pmi>�(�QJ�@�1��?��|���R��6J� �����	=ui�f��8h�jipG3��>N��<�R��k?ׇ�k0�?�l���+uB�"��M�Q����:;��E��
��!�kE��y��:L�Hm2*��R�~�ʅ�̙S�K��(��M�p�G�Fl��q�#P�^h.M5�j�Z��%8C��y��� �Zq(p�Z[W�^'�HHj��C'T�.}'��x����ء�	�[i~�\���7iO��p����*�?���{�a�_0K�,̬ջ����*�{��0����糁���]�$7Ë��(_��y�F��Y�PA{A�7�O�@y:�
fi�J7��_��BĄ�Ƕf��i�|����_��xX�m�Q�NO�MPp�3uV*�5���+��N�ǋ�f,��ms-�w�d�fpN�$�:�OaA���r/J� ���+�S`Ô0jܞ"�3T��熄��X�ڱc��=O��f��b\̪�:l�?V8O�r�N���E���;�AM�e�;��9Dw�cl��hrz5҅L>�ދ[���QŁ��-�nhH����ɎQ?�b��'ܥ֫$,&dG+�>����\�N`�Ō��t &�C���Ӊr0�c�8t�7-�A�����0Kq��z��W��dTw�rF�gJ��Ϡs'�6'�DG`�7i�s��I1�u����k��� �J�Q�Z��a;^gԓ��#������"�!y�?-E�W�;(��*�F�s\>-r �:��\y��#p�w��I�x��AV����w���T�� ��a��r���=�n��zp������bc��Cϣ�KSv���a�H)7���ͧ\Vm��9��%DT�cJqfG}�/���mΩ\�tTZ�L
�Ay��8�2�7Dp�{v�\dV����#s� �m3m"w�ڴ<��[��G�YF,Q�3�:�i�`�x~�
��c�^�&�P�0��=s�k�s�b.�kt�E����Z���:�o\[���:L�C�ަo��l-���[qNq~1�۾@Ҍ��:�f3,*P��6�L�8�~ģ����=k6��۝�8Z����J�P>��Q��	|F��C���?s0����q���K��*�����GT~�c�v�nm�LQkͿx�_��y�:-�����v����_�2����֖�QQ3��ā�?�ߐ�<��}k�\�q�g�D��ѥNb'������\L�/�$�O����ğ�Wn�#k{��O(����t(�?U�@8�iz��ޤ	�C�N	>ѵ� �Z��A�wcZ{~
x˞��3Z��e�U4�#:~dRf	�.�50D��r��5�$g�x��֠�H�������t�&&�I������4ʜ��,����.Ytj�
�b�@cZ�T6��c� ��[z��^{z�N:"��^%2�w5�H�8�ё�*�,ҼO;�ʪ�]���.�X��V)m($�o�AKCu�KE�48��N8<5��G���X����Y�����]lp$NH�����S�]�ŋβ��)��){m�HL3�};��v������V��60�o����C_κ[R{J3o���02��	������� ���YP��?\�Z���78p���M���9>���_j��쩥�,N�ܢ��A�^;��c�нR�3u��=j�Mz'iSi���L�D䰷U\$}̟��8i9��渼#)�T��Q���E�2�	Y$R�Y�_w�Yb�{�*��~��:�C��D���
>��������rf�ՠ@�&NS�2Gz������1����������B��JOve!�]{�o.�BV�/���5�j6,0�ٮ~�y(�1>�&ǟ{�%�Ru��N�ӎ���ǹM`�6{#�R��5l��$��3:@$�0���� tα�]����A�_I���ZPL�Yx�����Y}\L�	���q5ԗO���#\�l��|jjb+p��s�b���,���T�~Gp(�h�8ǁ���<�w'��FQ�j֐M�yKBo-��i��MgO���'�8KWB"��g�+���C�p������5�	�3;6�a1�Q��=��b��-�:\'�C\7�����ť�����xӆ�/�{�D���S0�l�ݺ)��ij%�n,��ؤd|t��yY͗��+�C̣҇0�q����w� ���;F���/�\��z�_5�'�뺄���C�eg���1�P̮�َ�^�_�7*Ugݴ�g��ޚ��UIZ�����=����s���8H�K8Űo�u�-ZQ����7�1!.�_KJ�}[A�h&���B`p�<��!m�0WV���	X)�b����7[��|�pgc��_�^��~��\B
���ӎY��⮗g)؍�|tu�@Z�0��_B��4�1�0_����#�:]�:���<ab)���)��tz�n>�� �'�B�Q_k����(��ޞ���R��W�ݫE]��҈�=�Bh�����$���/G`՚���=T�w�_6hq���Oۺw�%�!�^�ז!8�D��\)I��5û�sE�A��,i����oK$��lޕ>-�<�K�?z�a��U]l2�?�ĸݕ�޹�Ij��а��ȡ���9K�M���?i�$���mC�0]�����+r����D�O�vwd�{�"8&��*VE�֧KO�4b3pST��37���7�4�����C�4U	y/d�n}/����(��M�*��e<X򷈀^�X��~z��!}��/M
�J���
�g��1�&����	9���ڿ���M�vӧ��l��3��2�%����)��K	�%۽WG�Z�)<�-9�:Ƶ��ر1��Jd��:��vݫk��$�1(�U�1:)#�}P�����i�r8XM-"M��zeŕ�4�L���E�9q��[�iO)kܔ�f�}r�L��LT��2(W#�UA������3*~*��k�a��A�O=b��R ��eިDl���D�-�q}����rК@�}��F��ȲL�7��Ļ�]�i�eB��vWE>�D�����V��F���.�N����_�j�����Ū�#�c}�%2�9�B5�17ژ�+ ��yi������v�`ګ�\�zΟ�E�?Ίw� W�c����Hn�5�dA��f|���NK$�w[�����?��5f��Mp�<��M�������O@;x���N0���kp�v���H�V06��-M�$A9={<��X�ڇ�p�ZiWx�2����S������6S�pD�9b�f�^#@$NOshGy��6�f�N�U>`~�������Wc|bnT<����G�A C��݇� %�
