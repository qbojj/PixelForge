��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��g��C�$	��&�1�noX�j y�{���(�����:]�2 ��lY.�~wj`����T_��ڑJ��K=۞tN#1�B/N9����L�s�]"6HZOT��L�=��W�S�id�j��|��_�z����4j��9��=5P��<�_��4��~�jh�릂�	�-M����[ � �p�T��6p�
N���)�wT@����V|R�������e����n��_t�E�m���y�B�Zb�5r���v�10��ن��+U��������^qF�k����IGgw���*���,=��p�{_���]�3P���Ib5:̿�>�_|������(��݌��e{�&I��7���n9k��E��$���d�i�Tq7o��xM@<����_�ҩ��TcKs{�׳���y��ӭ�ETZ�Y�v�|X}���~_�e����z7S>��ŁK�eI�8�|)h�b�$r��6������^	���<�� �ڠ�����7s���	#13(⌾ؗ>��'�]P>b���_w��Z�k��E�i��L-��C�dk�����(�
4"���n(����*��Xz��ٯ�Q6�j��+��;Z��2Ʌ ��xK�nL�)b`��d�6=�Q�>4�י��y��) �W')O*��X��J?�&9Ƴ,�W@���H{�hx���D����oT�":�.e�e3H�,[>K�-j���^l��[7�^���"��*~=���x&Ƭ�2Ch�A|o�J�J� ����a8��:xxQ5�D�W�G� ��<o����Ϻu�g�K87vɊ\�b�Ɏ�������頖Q��NQ�}l�۩|�L�r�@��M�$Z)�MEEȰ�N�囈0���F�s|kB�q��aHloh�v��zߺJ!w�Y�j��W�
�S�gm����i����sCb9�V�[D�?cw����t�_�f	��8�'�#T�d�Ze�U���K����0�~����13�{��'�䮇��͡6�����yP����DPCeo�t/�4���\o+F�%.	D���������f�lK{������y��'�Mܗ�[	�����%��y��<���W�!5d����S�6���~VD �#7�~�c��A��W~6�V��U�'�B����#&�%���a�<��NE�K_|}���=��AѦ�pꆂ>%�p�-����d��\l*���a���g��ofᅨ�F�`��dw|2��y|n�)+T�>	}�404u`��b
w��Vd������;műk`� t�0ѽ0��c�)A��T$��0֎'�ܖ��u��XݢJI���u���1�/�8RU�3�?���<G�:*Tj��2��qU}���|�k�o�H
y�cTz*؏�ǎ;�����Gd<��MV�Sp�zg��k\��=�b�@A����Mb���qX���)`�&&��2e��`�edh6�U���Is�|�`���_�lc��%P�t�OD�д����~��p((��\p̍&��L瀛��?M����:����2��*�$��!�2:z���8󛌈��:bF��`���dM6�xV� � @/�HR{RJ�Y^��ݝӮ[��CQ�+V<���W�^Z~���)I�G1����#����X�d��7��9��&)@ ��Q�#��4<�]�C��(D�B�Z��su��
�<���hC�ڎ�L���&J���h�)*�9p	��K�H �	o�^���ڭ�D�k�;���^����,��A���ׇ]��dࡧ�G�	��q~z�E�i��/���
��Z�3w��Z`�#D�n�:$��搫���� �"f[�!P�M�/*)�6���M\�u�75���Qz�{A�w:�-G�(8��#o��\ږ�M�|	���i���cy�ȱc
T�i���Z4S�F#Ī�r��n9D!�������x.p���� �~�{�iz�Rg��.�r�4��}x�q'8�@�1�P��Fn�}��
u}(�y��A����%8sŒ��+iI�X���܅;4%n9�����Q�*�����	��L����P��E���l��d�x{�HNZ~ ��
��Hk���s�_�cH3�U]�#��3V}/��f�?ݳ�ipu�)F���Vx��<zɐ�P�����ʅS&�5�vi%ƽ���I�q�B�A��������t�9ԧ�͢Ƈ���MY%w*�כS�`��i��� ������z7�ԩ���k�`�ʨj�N+��SV�;���Qj;k�u}+�ԦI���a}Ts��j��q�,X������`��"v�8�]��R�Sz������N���֨�.S;��`�H�q㏭�B�o��`(�&���-���-���bz�q��};Sl��:�eR-�i�\�6��7���ik��7�'��I5������0��C�R�C�%Z8d����l�'��Q�y���I�18'C�+1iJ�1G�pW��۴"eQ�F�9�E{�81]IM<�B��$a�8rIA���>Ep1xt�{)�px�r�$�K�.�e�ݨ{q�v�ΐ���=FֆЅ4j�QF|r��M`ƭ�*���x �h�k�dw�8�^ܰ)�t�un�p�.N�/�6�����f�������Xv�\!f|�q��x��l�q�c���鸍���[�f�R��ؾ���S��U5�x`X�d��YRXa���P��ּ?��Ǭ�X��Y��m^�^��À�6�;b�����h�����cf�"�M�2)�녍]�����u D(���G|���e1�����읪�>��EMxx�����?}}��|��/i���F�-dovw��lBi;Kb�.2�	=��F5�ERyA1�I.����ۨ��)�7�t@r�r��V���V��C�f�f���(�)�Q��YI\E,�y6�'��c����i��5���SG}�[Vr)�v"p}�Y���0����w*P�'�K.!^)y�w%,�'�����
��8Ø5H��9�OD��s�y��@>�|�S�$��{�5�>��� �(~d?l�y���ǫ_&�=ܱ�p�W%-!z�=�c�o��"�[)��A,~k�C�;��j�]�V,q;��w&�E��9�j�T ���9��	^����
;�X��omX߁X�����i�+�t8Ks����E��b�m���j����7�Fp�c��`����ɭWc䓅���44N_��;�p��wh�:�fF�[
B��O[F(l׍�)���֡Նz�k� ��7s[^�/hO�2*b{?r6��~2�ڄi�U���֍ή�Ħ3���#W6�{(�w 7�x?"jZ}��A��7���}��������Mq��R@��_���򀆭&��
{ߦ}� ˲KG�f'�i��B��<���~A)��N������~�Y̋D��_E�S�{^�۫�r���� ���h˻�ϳ�R=�1�=���:m7��Mzq ��B5�%�� �V��ʊ@q�G@�~���LQ����"c�O&��g�ti����ꞔ8�WN�z=�u�8�V6`xrzVrA8�d����T�'�-��j��M�sQ`����N�������}��+e�u�)h�.-JX`���5L�A��䐲��I��MS�!JG�r}ç>L]�eA�\&@���#��/���$�˵���P��b��h�VB�f��Cl��3`�H�O�m�B�r
����i)$^R�`k�	Z�9���{�9��g=���mKm9��:�F����˿(YGUk��;j�Sk��b.�����B՝?/t��j�����5ָh��[e�K𓋮���C�	4�.閝
���o���M���Xl):�r���Ͳ���jv������m�����-[��t��p��PG!8Ȋ����2�`�-]���M�h���A���nAD*�@~�q�M$=���N�.`�ɶ�M Ы's���[6j�+�UԪ�>��w�����4N�e��p�����p<�\2p:��6��P�;�?��q��~y8e��'�D4*��R�����G5O���M��3�`�	bI,8����2��o?   +U��,����M�z��+<=.C��a]�ղ*��n��j��;H���c��?G�;�W����%��s���D��8��V x�^#��m����^�����[L���C� 6x�"������=����� ��k��N�uR��S0$$ .�ɜgK��V��9y��`�C��V���-�qV�P��;�f�Y�x��k,^a���Hy0% ;�/1~_Eop�W��6�g[<,�fu?�Xg���Cח8���Nk�Ua�������º�o��"\R"��������IT�(�`8؂tT��9f�,FὙ��Q��"_���0�w����`���@��]w�˛��)����Z	lq��,�>GV��I*+����~�2��
?N֐+Q�gL�G��O������Q$2a�T^<���<�O�e�����g�Ң2+����ce0#��x&��F�@����1����3y����9�vP�:�Z��,n���Oo��Ⱦ}�I��yư��vPV�Ɍ2sVc������H:y�n"i��`t��&0�~;�͒!Ѫ
S��ߺ΢����Or(15th��B�Ί���=��])�ps�G>�r1ǌ�`c�*��x�hxF? ���T�w�A̲��'���E�ܢ�Px��P(�fo�r,d?�g��Iya;�R,����n7�'S&��p�������Ҟ�|F��~7>|�y8��^�G�������ޞ���quՕBQs�g�K�W�<iy�r�h2f�Jц�:��׮7ٛ�-���^TZ�~\�#�<�2a��cF'���؍f|u�+t��ٞ�����+��(sN^k��z(l��(g[��4���1K�����Uͯ�y�=?�L]�ۂц�ݚ�~P]���J�]�>�t�=
.����;Q���G�3��P�җY��bNXHB}J�r�� _.��ܞK��'0.p��h�Hm�~tvT]%�ϝ��p&��������[����7�d/x.��E��DI1׳�+e�kFf6�{����hGC�Rc<*�J��_��c�ť<n�!�-���y_�34q�Y()p��8�h�*�t{C����@悌�Ng&�n��^���t`*
�j��-e����X1V�	6z���
T�1�3I�m�S�4� �{/@���'bTQ���p)��d�ߴ��{�h徕[�|'x� \FG���1A(I��;b�}à��N�4��ӚH���0j��^����~����)
�EI��E,"�͚_�Z��+��9���ZQ$���Z�?s�
H�5�-����W�6��~��v�x����M�lKU=��w}�Fp��h�6F�+0T��H/@���WM���a�y���s$�յ[�K������|V���ސ߷YU`ְ�лo����y�)�lohlwQo~��S�=0m�*��o|ރs�r��d)A�04�bo�	�>����ne���u���k�p�Va�#���8�Q��s��ˉ�kt���
���Č�FIJ#��`�����t�J<��b)Y_�{N,G���1-/�8ӎ{ߙ��j�f�R�B����ӥ��FR�,l�����
��|�Q�A�\\a�9��e!���a/qZH�=Qu�P��0���iQ�KVimy���g�+�;-���t8뫵+�$v���e��	hI�ܼ�h��?;-��[X�-�J/�����0����C���v��aZ�@���O���*��~%f�6�-ҶQ�WյLk�ƒ2\���i=�m܎e+K����rw�p�t����Tt�F#9����Kֳ�D�|�K�AMm8���_�c�+�]Nё����u/h>=��$%#�_����Ā	�_:�qJ�I�1�GN���l���ބ�-�I����ׯ�KG
"��K�}�=���A1��:��B���ְ�NY��t��P{de�������;4i������� �Hι�쎵U��+J�,��՘�;��!�7�É�l,l�����6H�#���@���+�B�F!\Mj@�,�*���D�-�ɺ��cE�e����](j�R,^��~���%4�)<���4����oM	~�PeDH}����K�р����=��gd�x]�? t�2��. �I�B���WŁ�Ko�+��}6�����c���t������e����-���>��1Y�[��)����M�v��_V�:�����w�V�
�;2׿hI�JHlQ3{̀,U���y���VsBqwf�������*�*�}%0#�}qcg���G�l�L{m�%U�����Y�r�Au�7.:�?#4���,ad1P� HȨ���Y�4ᖽ9����S����kl|�JeZ��3��ovcTG���U'{'���`uS�$��ު�Γ�6����*�ߚP:(���1Ԭ��&��"$|�g�i�s�%�/KFv�{IB�i��?��ʞ�╁rӎH�\��a-6[���x�2j�(#v��Ez
İ�0R��0}nG^�*r�UDl�88Q^��L�j0��p��Z`�g�.U��h�i�`uv3�3I�4��֤�����:pi���~�d�@�a��9jz�\�T�ovsƲ�%F��}�g%�a�H݂j�idΈ%[�9}�i���;�z�9�r�)e��s	�3F����A?iw�'��`��
j��b�9�!�ZB
M8��"�U���uUI��(��#Cj�&�G��0��pgW�G�\n��ڙ��vN�Z0��o,�l�&�U�
��|+˚g�ٌl�^�� �S��/�2���6*.S�F�6|��}�=#������1H���ݨ��yk&��?Y����V��V�qNs�Oʬ��^�Dy��	v<G��H��v��3�w ?����q���Mh�v�pO("�`7�\���I���ŗQ��r��Ӡ�SƔj�0���"X�'�l~M@����ߗ�9`��g`j�iwk��{�#�%�h p#�K>�O�nZ�9-E����m���USa
���~ ��JMQ�J�pP�f�;���y}:�)��ֺz�xm2<��ͯ_�I3��K8j-Ȉ�K#I��h7�>Bۮ���[��gY�p�_y� y��yV���I�4��n0ú��m�^��޾�s~�5�e�!�\�[��5������ǎ�P�]jpDk�OZc���WWUjD@7$٬�%:��eER�o��u��A�S@b�B�M�%�2�$�?�C#�K��2D�q]7i�;����5��x�=��:˵��sR���_ߋ7ø��~�#%~�k�θ�7�`I̽)}Q$s�*�KP+T�c� `l^�Pk�U2*Xa�"�}��3̑mfJ+���%��1���T�Z�C�g�c�:�K��s��Y�i��2��<��[3?�~�??FA��o�ĩ��8�����^�<�1�ۭ��[t��  }���M3D�:����r�/�9C?�� &��_�i�? 5S���/��*�^�D؅i'x9�v7����֏sk�h�H/���2N_ܠ���j?�l�Ӵс�I�g����]�o�&	��6W_J�l�0X���$t(��T�����]�a&2�GE�j�������D���Ӝ�g�D����.��#:��/=%�����,��I���;67�!� މ,B�F��z��"�K���V�k�.痫�er��dBś��B��oc~84����[�^�ͣM�{u���w�n���P`��"�Qc����w��o��z���Fm�'�se���w5�\�yw{��	Cٲ�H:oα�E�a�I9E��$�&>q5x���8"p��J���H �+<�'�E\���Sh�'����{]��{�w�����/M�S��eֻ��vׯh��{���T�^~q#�4�ks>��3QVmZV>��)h?��n�PE�=�3�)��l|R���X*:P\{��zH���W!��5�t&��5�P6WL�ↁ�qٰ��N?��!k���dlF@chϱ�6����dYi���&5�C[��@���#���?�
�%�u#oSd���K�s�jcΦu<u5�n�0d�F���uU<��k~Q����(��^�{�ߊ�V�v odć��E������N�{s��=�<Z& ������2Ӈ���R���I,8x��?]������D��̻��W5�3� �~�|O+.�e�����b�wӺ L��1��)�����+BT�|ٮ��\dۍ����(P��bk1nU���O-S⯶�k�q?��ɕ�o���V����ؼ�٧Xػ�%�p̀�#g�2p�<����>RO�SR[k�ܬi�%��s�Qtn<kQ�N%(���
Am&���3Zig���tX����JDb���aXy�#rL��{�A�OfK�gΌql!�c2z\oK:��
�Ƞ�Ԉ�)Y/�zfY�T.Z�i�R(���o�{s�-�a��|���2iH��Y����Ԝ'��9�Q%R�L���v%�	�z	���s��8���ǎ��h����fְ�j�&���;�d2t����R�AN>BtЇ��4C��$�?�|)S**���m
	VK��}Ʒ^'���Ql[fr�Ǔ��l�4���*V�_�_C�B��ũ�!��e��):��矄E�r$H�Oa��L_,Q�9�.z -��.���	��(m�b�F�{�����E5�D�@Q��yɹ��枟M�3di��:B��'˴b�SS8�
��N9bw��_Ϯ.�<e�{��D��j�Ğ�����9FAE�_��<�
�X��wt��Oȸ>���03��<`_8��"er�6���k���نz5�F��ad1�\j�)|(�؏��s�������Tw�#(�#
�`� ��062^�|(r����uy!l�#���0/2�JؘpVm-r�-��2���������(<pϯՎ��}�Y6�@���̦"p����������� �!t����E��j\��-�'�oq�vj�\m��Ǆ�me	t��{����B>�=|3N�3���߼��i��+���6S�s��(����=��CzP�T-=�t:���8�K�L��Gѱ��3�cJ�1����{�	�� �v���\�;���}��ݩ��� �ȵr 55F��?���RB^l&q��,�u$�H�����h2dV��~v�im���5�� 2�*R�f�v�!F����q�=ph��� ;��jO\�H�Ls���-ON[i��R}�:޸�OC(Uv�;����p0*�!��Ka�>mq�C���$iWz�
�Ѯ,�����\�Q�&�ewy��q^��2K��l�pS;��*����4�ruY�<r�ƞ���;�/�&諸x�mmU�f�m���G����U �:7�Fٺ��*���MҺ1J�A b���Zk#]��R�G����e�����v�"��$绩���꜆�������Dx�]�::��^��R�vh�CH�v
v�^��z�&�~�f"����Sʼ���Y��������a��'� �+�3����ә�)��j+ُWB��ן�z����+�^�_�f��I�Q;Ye`�=����(������l-&�d�x�#W�ny��W��c���U;��Y�9�F�C�Q/�OF�!9}�}:-{Ƨ��;[9|y}(�ٮ6�.'e��L]�#ȸ�hL<�QZ���q�(������){2u�$�}�Z]��%K+w�M5��"����y1��Y9�� �w�L窔})��7���5EV���ƭ�����s
S
�C��٭�N/���^] g|���%&���cg��w�ߔA{_���扚Nޱ�k<�2e����7�-@!�1�gF��Vf�<O�b�d�PF�nUD�4�����J�`� W��ز���g��	�mt~������5�N�ޭ�����(�f�T##�13�KA=�l�R��=�Ț�︁~�� ����LW��_��l}�c+(���i#X���E-ў��K��!���g?ͪ��F6�
�ńO�!hvK'w�	�����0?1�o���}:�%Z���*�%F�ʣ�KH��͑�	�G��L0M��~�KF]�X�}�ָ��V�e!�i��ܜ��'���5�B�)>궲�2kk��G��D+��y�'�3��0�2Ա}HnPt�γoOF�u��%���u�_]6FE��3����}��[�s�)����x`���k��)蠱��P>�Շ���^E�y����,��Ƥ�/�»R�D��GA�{�׷W�|ܼ=�E�?�zH�0b�NO#�;�UjOA�������91��$�kU��<U���Mo-��@�'�/�U.���K�d���,�#��>zUg2&K�׏ȵ�O�g d�;�b��I����Z�A#�^��±�b���4��O�(x�l�F�2�ٯ!^CJ���������BD>�
ꭞ^+?��YuΑ�l>@���	X)�-�+~"�E�`^e̾]c�Z��,w��=_�m����XB��b��'��b�K�� E`�[LS��"���D��D�����q�X1$��'b����'�Mv��T�ݕ���1�`�lN�-n_��D������7^>0ß��ΩtJ/�u�;�ݕ���m\glav�7��t���T�5,=���+��n(G�^�Ԋ^��uvl��HB�ܓ#m7����_���[�2G���(�x��7{q��A�_)�(sR������ ��.��P]�-���%&���"�d�}����L�!�(s�p�u���^�@>������Gj�&��}S�'ݤ�^�.���y+�F��$]%�D�3���;#�܉�+ �m92���j����K�qJ]#�iq.0�Sx������M����v���d�����#����3WWj����XFMz�>gx��덓�����"B�������=S��4dK�V1����MZ2	#�j>N9+��ƹ:9{�h��ѧ<�dWW��[��(3��,o�EXvN��s-0��frhe�n�s$�v"�?)�{#�l4`�3y5:>��^��(�����{k�x����#2���]�&�(?�%mR�O!!H�#A��QN�2�u$�/t��YDqe@ڜ;9[�ƖR���	;v�� N�0m�А�Φ���4-;��o�?r�����Vr �/���-�R'��N
�3���C�-�r�<��)?�N+����B�,�\������P ��C��;b8�-���ױQ�{	p��b���9�j�g���R/��oY���p�B��.'��?ʻ�ޚ\���O��y��Df�o_�?�]S3^s� ��l�y�=�0(kn�����h��0!�C����ڽ��S�k�(S���l#���ZI1啐� [f���)���i_�xN{�>�rw����X���R3K�W��*�T%X��� ̗H�[��ú��q���PG�]�KW۽ i���C%:!:�Q�۾EZ���y�R���^	�a3,��V��/��c�P݂X��Ȅ7CU�嵇�a�Ou^�9m�]��HFu¸3,�XSy�[�J<�C	�-�53����j���z�O���e�eH;%�hnץ ᅟ��E���%?|�ϫ��ڵ�T�w@=�-��照-���{��ZUa�~$�����^2:*|�u��%'��鲉��ל"�]8��ſ�bM�UV�'����埦7Gb�nO�z��d��|�����tVxJOW���U�[�<|{
��-q�869�s���������#� Q���]���0ѷl$	����~/?�C��7i�>�h���HD�ʻ#6����h�y3��e�BI�t'�e?��h8��`���"Gq��U�Lۢˑ/-��/��ٍl�S$�);X 8����E2F#�!�@>��Jp*D/�#��&�Ag\���V��ر�r uY����ӅR ;a�n�Sn�u #��v�
��W�w;�|�x�q��hR86G�(o�̗�=eEO��a�zؒ�T�6��J6\/�Y�W�@��q��5?����F!L�2��*� ��1�1��w.v�;�ֺ�r�]g)�{��?���JȂ�0�u�b鬅,-Ie��%����m�-Y�%��6����~VT���|�B�7��2|w�� _R��Ck|3� /� mw�[>�����2�,��m0}\�D��M��q���wX�*w"�|$ ��d�=���R������b�Z�	�SmKjK������'Ry�� B!L�NE�-%  Z���0�Y<�'?�%.��|jH�Y����Q�����.`ѡTof �^��S-���h��@����J���!d�eh�^�a�m��#BQeʀP��6�^�o��Y�{�jc<ė�~+����mF�M
��,��{�k@�J�� _��1���@�@�Pk�*Z���x}�݌�-����%x"Xowj�N-$	�ݪM"�Kl�5M�j
Ļ�*�+�_Ӹo�����A�Gh�0�1��&���9�_��N��&ł��7)dlE-N�kc�i��N�>a�r�I��w`W�c����5��݆#C��f�Csx��_��vU��'ʒ����`��Ă��Kz���{޴�sj�M�>�\Q�C>35��E<��uq���O���r�}��,�׺�3�����K��xt*�߷(�����[ѩ�:���qÃ]7���R��P�˃�7Nq��-��
��:�0�Z�t�/�z/ۂ��f�����$A867l�d�������U5���U]ڂbtC����(���k�sEs�u�&I��S"n�����,�l���ٶypظ�j��r���|�c϶h7��$|l�@�
v�e��0b�dP��?�|O�fe�u�uQ4�!u$"[�țRj_��R��Ý�z�A?2��}x�W�J��	���CP�?b���Y����m(M0IzhK+ ��T���,��^���A��g�OSRҗX)�~�M��h���\C�cr��UKr|�wg���Hx����LeD�;.������%R��C��Dsr��W2�U�M���&��)°v�;��񄜹"�����q��]��0��j/��}�jb���/��|���P���ع��m"��D��C�t9�I�q�e������S^ٙŝ�ˤ�	r��4�Zĳ�����o%�а3O<Krh`�� ��h�PBO�[�y^k�kx��Rv�J�{'f(7�v��A��������~ͽ�R:�c�`�|�����m�7)NU��D���x7�;+�3�na��ePBHa�E������qO�`E�%�F׋�:d43��9f?n~l^�M�ps��o�U� ��v��s_-�}6yF�#�@��HI�I_t���7��pJl�����w�;��\��J��������؅���̰ ����sl���ӿM	zj!I5���x9L%�y���x
Y�e��|�y4��+������&S����oV%j�>S�ܿ�i�f_��"�d�a[��F�Ĺ�?���6���m;ӖfY@Hۥ�*����b�^�w�/�UQD gQK�* Y0U"�B���;pPN'd�l ���]Đ�l9 ~ǒ	g7�W�cg�޳�{M�J �e��c�U)�aW�2��<US�2Hv#%S�n�Q�M���H�<��	�1�$�uaݹr5Y�߿�}���!r4�ی0ivB��K��PJ��Љ��7����'�K)iBu��Cj�+^�^�`I��S�z�ݔAλ��=��&��6o������tr�*�jj��k)�^$�X�Q��Y�;����W]R��:aBJ��cW`��׺GA��r'|�T?5�Z�)Ա�y�1�⾩H�ia��{�qM����]-�\@�g5��{#�%F�DD�v����	���К�mW@{��8"�' ̓tOu�j\��bi������Ϫ���&������&����8y8*�7�t�g?ѯq��s �iu���kH���&��� t�R�.�8���rrp&��]�׋;u'�?�d��73�}�X�����wI9��q ���9/��w%���i�w�b���M�b6b �KG�5z$�J����� fY5��yNBq��,�8��[7c&*)P�������"��K!���}���t�A�S�n}�1�ז��&��t��ǂ��[V,�{�ƝH��e�ή�,8��~�h���@�S �f%��L���j�Pcf$��d4S�~ѱnkG M֟3��<qޘ���낞
 @��<D*�-�	���j(#�����1�"Sc���	f�TG]lAZ��f�4�c��) �ʳ/$6(����N�)�}�u,�;��ӧ��>�V�
����4�\i�iIi{�c]/���ڸ�0&��� ��p�u�>�b�M��� �^)�V�ᗻ���fة�e�<h<�#�6�Ul��1�ڛ!x'�لM���[�"��Ój��R��&�W��yv�������%qcØ�r�AI#N"e�}qW�`6r~2H�Ǐ��~t��CU֥7n��~Zo�ߌ58��-���o���>q���Ni���J��y�jz�Bv��t6���n�Cs����U��6T^��"+������..�K4y���<�c�4�-�3�:z�Je�|H�s.�w�<��t�I&bQ����gb�L~1[4>��Y���R(.$*���D�Ց�� ���4�(�J���(ios�B"fO2 [��S3��nbgaw��h���ǆ7ͬ�+*�쀉ۛ�&��'�IT	�=��J�n���([q}<fTӞ��A�U�/OF%���]���_!��s�{�	%bwt�g3/j$�L��qn�4����m�ҙ6C۹ūg������J�-��{A�w7%��Z�$�4�q|�=�>E��/F��BdطBT�[���VH�mѸ
�#���z���uJ���Y�����?DX\6��y��W�}�ݩ��ۛԁO���Xb�n4J�A���Ы�z�Q���2=�M=f��"��:<�J4�<�{BUo
�����C}�=�Q�0d���6;�|W�������7�,���7zi;���"���U��4�`��.��dmœ�rփV_�/d��_q����+�+.���0��rUs+�m�����UY��6�*���#���
�0��p��04���[�0h�:�}���C��� ��҆Rfúd7�j��R�S��4"�'�,�0�I���/M�x��ځs{�)��x�FzQ%���/S v��`�E'ꕛ&�=!>9��`�=���� ��bťM��N'c�ͬ��3��૑W�+������GS��CЌn�S�p�B$2����Wĕ�Z�=�
[H�Xs>��9��ϖs�:[d���8����H���)1�~��2~�4bv�}��6Q���H���U8��Tt�c�x@����4k��z����K)	���&�X2��j��xX\�۪����U�T�7�4Y���ƾU�����T��;>�� ��i$Js��N"�|���>���3Ma��V&5��p�?���1g�*���ɿ�hkD(�5�%,��四$�M�/}�hzzcG:�����F�SP�<ӎ��΂���H�	��Z٤Ok ��o)���4�G-n�P�K�en�vM;e��	n��J�q��e�;�˨����V�T�	"���\�1�r�G�M���bw�C�3"�ǝ��L�9/޺a�2_�x0��S�;�v����J\x
[υ�
껷t|Tm�p�0n�XX�°���Vg+��\�JZ>Y{��o�S�w���_v!��;2�	/z�d������&�E�x�e�ht���ٙp��R�%����-�o�>'o�%v,J��(����.m�4��
Og�n�+hcpGx����؊M�Y	����N�T���V�j��{2���C7S�[3�֖�Q�I�����E���J��$�1�Ǔǈ}&J_�(/Z[�<��?X�S��!����o|����k�Y�2$H� �LJ�C03�!�D%��8��� m�Y&]B��U�]��e������k����?���Tf�.�Q��ή��ВІlN�o?��jAI�	BN�*n�% �sa:�V�#����4�l����7���b%�i섂���=���/#�H���%a?2�I˺mˋɡ�,����y���qO>����p��QQ��_E���v�f`$%�q�&U`*hm~AN�>?v��e�NA�[Y�w���[�*�v`�K���U@9͞Kb�AD���XZ^���!p4�6������.|�� �����T_��lA���t�����{��|2��Q\�Dw^k��,�z��(�:e�J,-���^���ã�Oz 9���w�3��0��5�U��ے�+��!���g7ѱӷ�J
��Uu�[�l,��F?���1���LoD�=��c+�t���������o��HJ��O+�������۶�A���pO�q�K}Q�[>C����%p��T��� ����K�_/q�R���p������[�T���(���;\ ?�X�K�Ӏ}N��	���n��T[��^���W�� R�J� ��\,���1��ppĹñ'(LR���T�$�_짰�wlv/�9}R�����Bg��N�h���g����ތ�v�zs���Dj���Κ0_F���ր��t8�M���ځ�%����3�o��l0���х��������ѝ�ƒ�)���.�$�ơ�	���9�4<�=#���8��Rw��J����� �[3gm��O�TS���hVv���[����ɝ4�e@^3��S귨��i���=*]����<�\CԘ������VN<�Йi��l b�.%��W��X�Bi[H
��o�P]7y�ܓ���W�BF�x�_�APY�>�H��)�G̍�u����|͔�N���8;fF��:u�J/�Uws�Z/�o�wPЯD6�$�k�����t��;�Ϗ�a]�hi��oot�n�lf6>8m/����E5��+>�
�O�1�y�Zy�����$n�A�(��j�bĲ��𒕮!)�Ԫ�$�o���r`?ƂtV�vu��lC�3�ǎ'x�wu�>��B5]���ΰk���dو�37T��>���6恇�t�۾��1�����ik�F��A���M_ fcH�v�Qf4ؿ�����?�V�`���ߔ�8���U�2N�9�9$��:�Da G/���j)3&xV����l7st�*F}�D}R;FR��������S#V2��C�w�{V�P�e�W��uΉ��i���j��,�vyx#*�r�ihy�-��PtS���
]> )�>�]���,8�ՎΏt�`��[X�w�;�ݼ^���7����҂/w�ؙKN3��N�5�����U��vz!�,R�B6@H*^*��Y���Y��i��9s�+�*��x�Y�=��Nj!��3��.�(sェFM�Ϋ�&j���*3G=�d���- �	��	�̤�^Go�h���J��hٛ�Rz��4�ʄo�����`w�XY"+�)<9�@�0��6n0o����!7�FB�Cč�J�g�5�u(܀M�I��#����\7]n�( w�e���Ml�q���&��0�S��i|���L����Ŵg�C6�ߥ5ֺ�H�J�3�풡���M�L����pS��(ܔ��D����f2??��8ȢS3��^:n@^�Z//y�hVH:!�����E9m�Z׾p��3�c��� �]!�⻛�l,S�AY��EToGֺ���F� N�����?�P�����]�e"���?�Ǚ��O��V30�BoC���^eg�"{Fh�Ⲩ�k�SL�����~s]���f*�%=�R'z����`R�|�v�WOQ�T�Z�g	�qq���l)1.� ���͝H��޾�N�-���z�1�0gi�:]�Z�@�O[��n�!qd�ٻ�o'�[� m�i5��r460][����i�l%]���t��tSAh+��}|�]S���>�KE��&�Z+?n{��5��D�ɔ�sO�,�~)��r� `[�
b�i
�l��j��!U ����wE��<z�`�,>/��o+�3�~��1��%�o������ų�1m�˕��#L�tkЇzd�p�>iڛ��n�7d!>��\�p9"\$O�Q���#=*����C�3�~��Iy��2$����s�ζ4���X���C�Ӳ�y��Ta���S�yN�o�_�&KG0���X�Z�F�Ď(ܼ!-��L� ~��5ק�pZ#^!�[��&���'E���g�T��#SНé�?���I8A^���៶���i����J�� �?<�H�����ɽ{]T����5�բ����mRG3�}�3����A�*��oCحPB;5삯P7��Z5�^�3�,C��-�!�5�7d1���#���P�1�1ɶԝ�����+��''�(���o�Xm;����-�G<
�p�T9��M%3=QV�QC��>��8���,
�8�%-7n�0�V/�GV��CM�nz�� ����!�ZrgR,���&MÉN�K/�7'k�h_�ڐ�/~�ƕ�zj��o��(2� ��
���
����(�i����dy�e�}r�Zp3�w��n�I��Ξ�^���yp�>w4Hl9� +|�m�OЋ"n�_�[w�S]�zp MH1��m$�:�ߜ�5�+GR��e��>��?>�l�Ա�O�8,�,/e�`ݐ�8~� wT���y��N\Q19�}�;��DV3sKt��{��yy�uYQ�����(m���D���t��p��|���`���I��͹
2r��PaH���M<wM��9@���b�4x����ؼP��g)~W�Q��k�.��Ա.��E��Ʀ�fz}l���%@v�����2��o�N_��tH)�a\�r�p	QE
mR�*�3+;�w�&,&�9
;{���	j�1�$Z/4��-GQ/Qк�,R���J�����|�MfRRj�RZ���	��4�l��?8
��䒋%,�Ҽ�#�n\���Q���cB�ij�೼7�Y����`���E�.��b�PG:�w�y@nDOcIөʼ��t�ރC�*�ɭ�0��:J 9HX]F0�J��+��bAi�)�J�Oj���6#�F�M�\���h���(n:��Z��3�pJ�b���k����G\\$���:F���HU�3�4����#ʔFn~�;�L�Ҫ���G,
�N�ni��#c�"�ʥ����4 ��K"�V;�g l���P=�|FB�]!��sLꝙ�Ig��Z�'���:�)M��?�HKÊ��#B����
�WY�#���Սo0W�[�� �;>�K|�4�s�î�z_WHUT�Τ}T@
���|�&Oh�7=聾�B��$(��tp1Q�����Sp��ʋ�ϝ2��o�?}X��3'�;��KZ���R��woz�mRO�� �vbmJ�]�+��[�2K�|�h�}�SD�'H��&�;�Ax+z�o-������K�<�jJB�?Pa	�l�Ͼ �R���@�P��/ �Z��:+����=T":�:��^������n���A̒b�������H�Z�%N"����{q?��\��H9��sU�n����l�N�~0�J������6S�W�ϦV���5�,�ڲE��:��9PX����}RpN���_c��c[��OL���Q5x��KS�(Bߌ����t;t+�������d�Ry�s4��e�r0�����|=ۧ�E�n�4�(�!}���B��mpܓ�c���s�D��D���x��vN��KND����G��T���ƚ�G���VE����ld]��k�������s�u��Fg��ȅ�z��ٮ�c���K�+nU��qE�.�#�̔(����_����b���7S���5w9����M��Y���Fv�����5�Atv1�|�˶�sH�=s�BH���.ܝ<Ko^�-uqĝ� *eEohy��n�J_qL��2	��m���*�}95 q-7FJ�R�=g��S���[-=ޢ�V������Q�ǟ�/��EaR���9�$i�l-`���28�E��4��(�w���hT$���V�:7���[$�98� �b��J�h(yL��uN������K�
� Q�/��l�@�����~���`H���O��	k���-�<Ś<�"S#O��ܩ������f��\��1B�O�%���!`�����j�x�x���N�E�A���\.�S�r"���B��\��Y�cGj��]���p"F<o���h��o2*���p5�^��n`Ï� pZ�ZJ\%C�4= ����0!��j�Q¬����<��_VP�5 ���q4�u3$��=����qI1���q?!��e�/�֫������ +O��_opX�_�U��}���"��M1z�������t;>��K���LR�٤ ���V���]ŊPd��Eh龕S$��^���-�^��S��5;�+����6�T����G�)�7�L��?���q%B�5v�2,� o�����,�,�j�`Qa�m��'�V��Y�����"v��avxo��:����
����	f|&�D�$������ �)���NR��\��_�r7D�K8�|L--R��9��Z%KJRZX��$c��?p�etc��9�� n���	��\�m�ib����y�l�asm�R&�V]RJ�`��-i��JM��k���I�����%�Wq��K�j�-���B 3�f���G�p���b?̷���z���E���Ӕ5S�,,��
r�WC����^�2�y|���+����K����O��߆N������Gl�ذ�U�W*l����,�=~U��I�R��;=Լ*3�Kbk�>�2�'�����̵���Yz�F�Z!R���5f�@]P�,_���b:���
��� �XaU��)��$�����%ؑcl��Iʅ
��iԽ�����B���3"ĵhw�H���<3��Ƥ�?O~��"���sR4YF�'e6��Fs�6����U�R�<8��[,��N�wx��3������Y��c�0G������4�{���� i}��]����j�ᶂj��4�rҥyۑ2��~e��p|�j��'Mͷ�^��c����V�/8J����T�Sz���9.� �y�Am��Ҟ/��C�P�)�
�H�v���D�WU��M��.=�WW��l=��z] A�\LٕJs�x�Ґӕk�?�?�Fw-���9Rj�5 .�ho�|r�_yVHF���P ����2�'��������!���}�-Ir�j�ub����m�!X���!���$�B_.��,�<#A�E$�S`!���Xj���`T&��� ���E�VPD&�*M�%;hĐ]���vf��ϩ��>�����1B�q�e�%��oR�)��8�e�)��l�dH_����V����nV��� *� D��$ڟ�
�����F�6∭���a�`�ܠε��MW!q���+���޳^H�η���SU
�n�=�BkS�F)([�_�m����"�{�G���ׇaW��9dIUY���7d8�[�b�ugZ�aZ���v=�2�����ȗ3pf�J�3����L�Uם
����?��"!�]�e��<��U��'Y ���]�q *U!Z�/3&�]��7����6mKP���Xع;[���S�G�ً���A�L/�����)�:���	Z�i���g���F�hA����n�CB�<��/�d���)���Q��Rh��-t�2������ Op�UK�Z�_��X	��ʚ���,�&��V�K��og�D )�cC��Ɖ܎Ge,�E3֤��ƠY6H����|���6i��V�yo�h�Uи<�Ԑ����%\��R�@7���fVs��7=þ���Ǥ���~�{�̎�y��?�Ĝ��gE&Dt�`�kWm9a�]��r�	 ���^�����4�ѕͲ��r����D�rG��9(ޚL狀V��3���˩��E^����FboW꿰s�M���-b��+Y�H����?�䫖�*���P�mV��
�u�b�N}�������
isO��L�		�Gɸ{�	��\��]�		j�˃W���;O#��\�K�Y7�6Sk%�#�v���t�@4 ���a��F�6'�6a��|�M�1�#��mw=wC�+n=m���:����s$����L[SzB�V�+{���5ٵ��jX�zcJu�D�	e�w4���%�ڿ���3�VB��� #�'L����ڃ��s�e����ƇpN�������@�}���Rd4��|ggz�r������a_S��0li�M�w�F�F����� ����ڌ`�C�r���J?;��6x��E�%������0x�N���)��_�c�2�,#�U�F~�}�����OPV���3\��M�3�1s�%��C��Th�:�7@���rL�9����7�b�:8˙�������4�(���1y`͆�$������'�\p�jM���(�,�w�je�>�f��������uď�0rM��k)�_m�`���4����Wa�'gCȭ�&�s���t� �vw @����'�Q����Ϧm�ϫEQ5F0�J�g�,�M
��Bv���mƜ�nFN���ġ�h�`)-���"8�-�� �u|&�b����2�N����RW��b9C:�
�?�_�	p��O�{�9>̪0��i?���q���k����,m�_E��,d�t��g��̢	�*\jd���"Mp'��4O+wc<��)>�e�AA�@�h.��=�.Y���*ͨwf��^��Q�V�;���D�Ո ��!��	&��V�ZJ��$��N?�6-cdW�j�E������8|�k�3��Σ���N%�(�41�ɰ/A����Ш8e@�I�!���\������"�ڳ�+���'��3�JmD8"C_��A��}C������<��^	5��J��b��K��pN(�2�e�.�Pt����ieb��*G$|P˥�_fP���!�8Z`$/�۷+]ñc��De�el�#&4IГ&��a�ފq��1t��ہ՞Pޢ�U��������{$�^���::�rHK�	���$�������v�K���b�6��/�>�z�|~����䕘�%���=H���;���]NJ�L��sY�xYcs�&$B�<+_�L->��C���py-�7.��.E˷�� �t�~gn�L5�Agą�����)���Ęo?H$3�_���'K$y�W�m�RzY�h#�����Td8� x?��x)אA�o��M@��ك(�����n���w��	���9N�;�-���lz�EL�w��o�0K���� 涋�j9��� E�!w<����+p&��J�eI�Zҩ��ϟ��I��/
��4�q�@h����:�
���S��V;�u��jX�s)[�,��5ۗ).Gܤ�U����|g��.�������T�E��7>�+W*�u�$�cg�p��E�.�E�e�,b��Yw3�$v���� B�闾���]4��#|��sҲ��dlu��Au�3�+iP���|��[�a�1jO!�1�N�U�?^G��G}X�P�t(��HQGɨ�K����A�N��&)�T���r�>=[�da��~)̢�1�����F��7�ߤ$��\������|�v(��8xgv�T�u��\���j��?Tçf��1���ȸ���TZ�bt��h��]�&膾O�`W~KU�S!֟Asz����{W'�!�-�����R9��V�`����%��Ӝ��V�u�in3Y6�("�+y��κ�jX�'��v:	m|*8�PI��~w�}�f�L2���u���B�Ͻ.��}�L8���	�Cu�j�V��L[(��Ѥ
:�f�6���,'B�X{:꣛�*a�g������Fx��łՓ�e�[�y����:"O9��WJ�z$�X�3�Y��X��i	��RU�"����jn�� ��..�7>�j��N��OA���d�x�;BL0�Ĩ}�qB*�$�$
�~�� @p#[y�emenZ�ʺ`%O�on
zX&��(�zT��\�kA�A��xt�=V�d��$y1�u��Vr�.���;ޜ4��Q�fUh�7~~�,��]d&�!(�Aݿ��ӗ�T���6az�lY��F�*��/଎�c�a��!A�/��ڃþs��R�+�w���Y[��(�b�^�s�Y�_�Ξ �����@ӈ��?�T��@+�@_v�Y¾\?����xZ�'��ۃ*U��W�
�i�ٻe8��;x/4�vW���-����Y�M����#f(��O%�s�7Ǹ������aHQ��ta?�J������y�@��Y2�A�z�!g�F�UN��pYYRR(��8�#�O�z�ll��8�)e�E/?�'�:e���Xc ��|�����'�Ҝ���WmDgy� �Ż��lV�n����)(�՝��d��;	b��-�r���/]�|�A+��d˼��[��Fւe�6�P6պ�~�p답�M+\Ȳ�ө��ܢBQ;��@-����8^.$5����[�^�O�[h�ɯ.���yW�}�3J^�6�G,9��8�.���$�7�g��˙6���������ey�&�MX�/j���~��Á*�t*���8����9ڿ�R�Sh=��C��	yJ��Y®���bߧk�x���ǖ�%�w���"�����
ބT�s&��.��]i�$�AT\l�F��n�cmWL���.�U��ۓ�Vj��o�{��S왃�H�3	FE�#�αeP�J(֚h;�����[��B-"vq2OU��|M\��ʢ�l����yO��A�P��'!R�?�HH��+/��oއj�"^� ��ӌ��L���\Ɵ�5�'#�d1u3
ϲ�&
~/�����/�%
GB#��,�7�5��u���.R��/b�� *��Ӎ��H�d`�<��Y�+y�����#�br/�����4��t��S��h�_�$&�:BD̸��} .E�Y67=OL`@��S����7R��Z�Z�n敔V��q�
q��m,Dn�ʢ�L��7�X�5�j�=4����@33S�(؏i��sD�����f��� �Z�ǘK�f �c�<����E��L	��Եs��:�����ϻ>���kP��:�ͤ�)NXV�y�+l�p^��oa{1u��6ToK7p-�r ��ֻx�zϵ����������m�ɬ������W�VlۣIn�Y���M�Ml\�tR)����p�$�<2�E�ϳv,�a�;�~�	ۊ�gz;`�(,��ʢ���	�x��.΄j�B/�j����3w�GX�Z��m�q�*.�fk��~0-������>2|��3�h0�:�`�\�P�J��h>�,w����}Y�5�`�]M�V�1C��I�TB��zB���D3ᾉJ3X�Ĝ?cޅzH��܉3�0�5����V�T����������i��J�϶��I��ٹ�kC�uP�������:.Ʈv8N�gM|��
� 3%(+r}v,ݔ;[!��Yt+&	����\:F$d�IJ&���2��Ks�G�� ��*|>�Ց%R�3C{�E0}k�(��K�v1O˄z3aBzc�����\�ez��H�j{�?9ej�>����A+'�A��I7�_�.�3G�Y0�5P�K���m��z�)�Tq��FO�i'Я�!�s˗�R�N���Ѷ����!a�1&�C�դ����a�{�P-���J��wq0}p-�CfҡZ߿�V�1y�V�7�p�Z��qC�͌(��ĳ��m�W���X�,.�N��
Q�7v�������݊�zIX(�N��]��s���aNZ���f���7a����2�hϝ�k���WRC
)=ʡ	��
���Q��s����F�4/����7p�i�����=���IV#�>�~�c�MJ��(f�S^��j��T5ho)+�1�ck QbY�G�@�M���G��9%�D��C��[�׈o�U�4n|�����R���J����Ex���Y�f<�������_�[bP���J�j�o	�9����ѱJ�� �__����:���B���V �x�aM��R���7M�$��� !�%�!÷�Y����'����$��^;���s�D�~OPk݊������C��w��k���~	RWk���K�}�\zƆ$����ɘ�&&)�Q8m�!����u{�̳|�*Y��D�\�׻�2d��JG.?��M��3kˁ�CTlVY8�!��[��s����s3��U�੆�.����0��c̞CKR�՝����ծ�<���_
w������揙�3��&=B�yM��R~���n�� *�e}lv�G1��w�3~Cઈ�ǉ���.U��e�{�c�3���� ��:�9�A��9J��J��C�@G/�ֿ�o1��j~-��K^]So�`сTq�K�ƚ;
y�F'�G\:P�S�'�J�#�>��|��_�+�$�����A���JU��ģɳ
�tBa���nMxu��6U�j���uh�n.�g�ukIǻ@X2�3�����(��/����i�^}�f
��M.+�u�>J+��7��1_�:3��w�� i����uk6���ٵ珽�xRՔ�@�Tk�j �aQ*fM*i�4�M/�Dw{V5Y�S����f7GW1������(�^�E��^�9�B��o�K��	8{�����b���JO��İNe�:JɎ���a�zlXU�}+����i�ڽ�x���HUͻ������G�&V{պEN��-ֹ\8e����Z��!��v�	Z�C~�:у4<�z��R�cR��*U��bje�g7�{>�[�t�	Ŀ,\��Ч���j�	s��yi��`�|�3j�~��M1d�@VnÞ�������Յ*�֠�9,���@�ar�hF�5'�˸�L�7����?�=��l|{������qsČcBD�w��z D&p������?~��C	������#g`�a�K���k�D#��z*��]aI�	[t��τ0��X�aB��� y�'7��`G�Q���L���_�g����L5�=�]�-U����$0�Q��b�I8�f}<�&�����X�"=���[!������;5wм�DV�­���VX'����D����DACW�� l��q*�թ�Xq|�:��,7��Ϗ���_hf��i>��&��H�r��o���e��<�UO��!m�������@3����^�)����췼~��&�������)��`�*�g����>mqΖ��e��uc������yntf�d�l�+E�b��*��['�J���_���P�/��~J f�Fx�0�� �� �C��n�!�>ӇΨ�h="LnhEEi��K�O@��1�������g�8u���|�z�כ��P� ���#��p7K�-����ȃ<�up�?Ւ=W��yE�����]B��k�(21@�gs��w9��HX-�r�x�R/%�����d�R4G/G��=QK.��k�!��}�|HW��IyZ9��R�������	��O��#-r��)+�����y
^���TqR���N������vNޥ�?���ި������q"<50�]�}��ޅ���@fV30ū�E`M�MU�q���j��A�g��jq5t��suA7�ـv�
0I���-
�B��RR��P�?��؀�N��u�xϼ������1=;�6�a,)�&�5'�X�[�5�b�&�A�\�Z0�����t��^U���}��4T�6��l����.�7(�*[{2>/YGa	)�j�,#\����5�_���O�<N�uC��L`�q�#�AW"�/���Oh���� &��R���Q���YCrP@�(%�uiL�aH%QI��~�k�f�!����W͍N��8ͱ����������q�A���J��h��ƕxŖk��@�n�`�ބwu��{̜�8ϯB`8�{§�hWU�UA�
Ѡ�����I�u k0>l������Ӳ�Aj���|��-c�=Ų:[0=��®��/}��@�b�����3�\djT�P>O�dC�U���ֻ��J�C�f޽E����q)�N�u�#'7z�	[��FS�ϠYm4���#n^��n㏾��BCh!�t��J^��g�2:R�[M]e�!ϕ
8 !�#�����V�;Bك*8�V k2�r<4��@���s������%��gQv�}����8��,x8�J؊Y`w'@�ڑ�u#<V("2�7��[u��r��l���oh�|b����m�*]��ſ�/�u���DX������3 "�t6�^u-k�;�ׯ��hܬ�+�ܯ��{<���֬�ms~����h�"IUZ&��,kfk1V��}�F���!�J��.�b8lN�a#4�ˉ��p~��6vG#�:Fg��g����^)0�?IF��A(I%�wF�u���C��o=3 _�u�3=
��8jgB!)A�����**P���]+EN�1�1�崝�Sh�܏9��gD	R�3�eĢB`�M��L_��������v�ѩ��RՕou�A��L�Yx��n�hç�g ��d�p�p�cZ�<q��60�5��)����MS��np9��+�H��q���,v(�z^󁔎�1�N
RE��ʞ���[A�;����S6�A�al�i�au��pz����0�H1Ex�7����眛�q�����/>[2:��L��\*�kb�����j��X�iB��r]�k
*��8j�����f�3�$)�N�p��������p���o�H��cP�d"�pU}CT[DD�"�SFf"Rk[ۻB5ڴ�5��R!E�������}�ܟ��>Y�ǯj����?�R
��^�s��zO�3{<MHS����x��c���"3=�$��_�Z�N�k��S��;7���.��mp�́�15����{�r��)Q�.���S���8i�E��GT̞����縜`�
X�@�|�t��)�_qh[�fK���?'���un�����(X��,�o�A3׻�w�3�$zP�@��6D�ʐ��f��l��V�e4��$�q@L|�j�Y6��S6P��+)�=!��e��-���ϒ�J!	�]�E����WHx�����X�F0�m`�_���
m��E�kn�"$��7�
��� ���f�!��Ō�GE+V4����-�{�\ 0�f2��t��ʌ"��^-�]hhI�W�kk#��@'��2S�8&/���	�	�`MMۘw9p���n����1
�2)lz��{-�f��"���j:�m�w@ ���n24�"�k�����>������������2 )clt��3T(.��7��E���Vo%d좺���,YR4N*m�� ~܎��;�-�&��|>���Ujb��:mޡ�� �;�M\%���d�[�[��Q�7eD�9f_{p3]�c#�����r��2F���X�/�M�t�JJ��#��S��G�}���G�]�8���*%�b��7HM�T< �΄[�f�1F/}�W�`ɤ=a�慀b��=��Q
�i��l�!��t�ؔ�3P}.c�� n�6aS���~iE���M
]Pz��Q��W0�U/UM�b��q�sW�h܊x���?d�24�I��9��K�����g>�/�&��y!�)1����F�4/f�/_z����K51�;��o����ѷ��5��o�v��X��ApQ3uu����Z��ڼ��}`O��
 g'3*�Ʋ�ё����y~V&1R��k����K�����x��"_��&�!���A}Z��j��Xj�&��b�/y����BלP"�M�8�g�<"Q �0X�t��3o��vn�_�Fi�u�������6 ��m��4���$�rp�H�XP������uTFR�E�Wg�;ẘ^��:�CE$��F���9W)� ,(6���:��Y�vQ��#t���k��Q���1cj�(2W�������z�S˹�5��2�d��Xȼ�&���X��ǁ�ո$O���m�H��	G���rQ�r�ɦ�Ђ��R�%�f(�e'�+=�ۗB����&�/E�>�ʵ�eF��pN�XJ��7JS?u9�7�M�Io��~	��wԤ��v�-��wܟ�*�F��Y.�������]z���L:���r-tn�Ks��3�F�&�_��{y�׿7٨�(���<U)vk��ތl��C�TːΣF����t�|KFC�����>���yЍ�2�ˎ�Z|0����m�M���q��Q�7�f�C�%Nn�,�}4�J�1rCX�2ԨګOv�~��˥ϚA��TAm$�Z�GV� 6%�PJЯ����;��1�k"ؚ�"��W#�E�d�!ρ真5Wr�hY��V3j�i���]Ƚ8ODI02�}A��x ~AL��UeI���JJ�w�v�(�g]y�����lʁ�.���5P�F�s��\����sT}9�)��f-�B����;��V��9vS������1�O�0����UB���X ��lH{x����le-����Zc�$�pf��C�V��`|�$���=���k&�J��C�����0��8�)"!^()a���mg���j�SN`��.:n����x�Vƻ���T`$m-������H�XXH�z޸\�*�Q�A��@�x/@�"Vҿ( ��k,�ͥv2�KH2O�yd��+�(�.����M����g��i�n� !�	��4� �ꛁ��c}p�܈e���{l��V�t�!/�
��Ո�d������m@x~"��-d)��M'$�z�X�w!zj�6C�H�5}�&`�˼[��vJ��4V
q9\aj�X"r��7���	��?.Zs�þ��&�eu7�
S'�"��yG����1������]y�"� ��+k|{ő/ǒF4A��^c�D���gC�Q�l ��&���nn���S! -���O��VTz���.la��}��Sp�>�Y����%�i�1~R��/G��������4ϲ����+n/eI����u�,qL�4�R义E\���!���|��䑳u����&G����4u'2]�[CC�^� DC�o���6
�����/�=�T�T�����p�VqX&���~�i���b�*�{�_��^�ܺ�|����t#��+����䝽=a*�ե�|[z������C�Ů�`!��+��-�H���R�$w�(5�;x�&+L�`a��+����^�P�ۜ�N��u�������K���n���1$~Y�Ĭ�\0Q�'sY�2
Y`���ZCT�.v�Z�2(D��Ojg�b<�֯�C}�\}_���=���c�U0���	����'�#�	dW]nb�\���I!!�K�߸o��c�bd=e[��T��Z�����гe����|�����+qwɔ�js����Q#&�j�(��ts+C<�[x�!���.<zB@��W��!F�WIt�u�Жܢ�Uz���[�00TJ��� �pa��;د���>���NlF
�$:����{kL϶�x}w	j��br�_3���ڹ�.(4i��p�h`Sm�<��5n��{���ٽ��u�c��̄�Bb�ڽ���ֵq%��/�`1�&:8�xޤ㢂�=}o��	Za�H��ߜ?*`'��q ����=Mטi=q�T����#~�ˇP�
�̣8��䣍&�N��d���Wʌ� ͢��̅�;�̓��1:�?�����vKfc��ة2��Rw�}��Ϧ�d�2ݺ�8��#jP�R�v���B]�WV�����,�`yc�~@o+σ�?ǈ��A
!��t�%�����bO*
Qc���7BqFA�����

��!"�x�8�Ar����u�m�������ːG�B6� �H��Q��\��P߈J`
���Km�v:I �����?�k���,��I��]v�'R��A�H���|��=k�ae1����@s���8pJ+��q:���%�f���/��W#����j�p�w?��d��"qX�@C�x���3��y7�<��� ��X�Ҵ�^{9�s��W{�؇�N�;\� �j�C���9Ӱ�A�{P�Q�øV]��x~ �i�0&��uz�m�m0ʬ�r���X����R>���C��"c�:���8@C�l�j���&Uʃ�Ї�5�q�aXZ���F|𡲽)S���vݟ&�פ��Q�{��gN�#�����	D�x���٨��/�5@ � �ߜ]�H~�D�hS ���|�󤒴�^Xv 	[��ˍk|���Ar��YǴ3o;چ��~�jf��,Ȍ�v�������6b�omt�b�/sv��R�&��=*4oQ,�N)%�h:��0�7�V����[m���?���e��Z(���Z�B��s����m�e��L2�	X~bL�?f�U�p	6���<c>ǫ�I����"�թ v/G;?���{��K���>�Y�b!!�Hw۔ ����9ft�r3����
�A�u#/J�\�O�֚��=�8!թ��o����ޮ�ڮ��%3y7  �nf�p��[O��ˇ˞���h�<4ۻ�f* y5�'�4�5�*��*���{?C{������f��l�R�����/��OcD��� �Z�m�7h<W�[�XO��*�OE�W�92��:Oo��=���m�� zM��u_F�=���V���I�E+p�m���p���,U�#n�1e4�R���km��K�����n��A�O~������(���FJ[�d��ԇ�	�A�.����Xoo����1�/�>V7o�}�V�7��9��S�i
��:*/���^���Ƒg)��e�?�@��q>#�;����}A���%�g��Fɿhz?�����h��O[�R�q`�3����B��|��E�G#���o���?8�0�<�,E�GXyv��Nq����6�9�?�KU�#hz���/��?Yn�C��_h�,.����9�hv_��BM�Z�j"����_��, =8�MJ����/�)��!V�cI�� ��|���F>� �V~5�0�m��v��ۣ�t]H�����*�Z%n�a���"����w���>
f �	Rp{R� 5�ΐ��}���r��W洑��ܙ+1lq��!���z+�����GD�#�?Yَ]F/l��N'���y���y�Ȍ!�A���S�80!K�Vo<H�A��e=�/�����ᒙ�����x?^Lx1�[��Hv�yH�[���Zt��e�4�|�X��_��)�T�hV�v�ƣU��g��I���г@3оFU')����U��7P(+�e�*s�Z�a��p��a8��P�}h��"t�栊�
0�U�#R��\>j����F���0�P,͞|���T�f�)�f?��㐱������8$���G��������K��m�n֤�ķ������x��J�`��"E!�����e{1a�Y�bk�-|�Wΰо̏�����Y�nRݧ���CM@l�d �C���!~-��H��xL�5�x���]W&��4ǡ)[��y���{�Fz�i@��)n[�5�U�F���~�m�1sw����<Y��1��a��qU.�����Μ�H#��.�sw���$MFX�}�r��KwT���t�v=֢F��5/�㡈�>>JjDJ�����3���*�~7-�VT�zS�+�@��L�̟�����=�Ս��s�}7|S.3��io��u@��kEK<�C6,��������B���oB��]S6�I�=2�,�K�����u��`�IF��I������M�H �(�U<�u�'����Ii�?)�?�����q�آ�zZ?�(u�v����}��ʷYΧ�`�Ϡ"���ԙ���K��.�-I-'��
OUR���m
��X������xD�&=�y���I
$�bX|���i�屝��'*ŎL���k�l$gO�h1'h�]��m�v:鉭��Z��6s]+�u�:p�A�B�����&~��Xbb?��x�(�qr�z�(���)dv�w,TȬ��S�֭�����A)Zm�Hq�۞���t_}"�.�E@�p���~X�*�q��w�mN�3<5�T��o�q�D��:�z�_�kQ	���X�.H��~z�� �~_�R}����"��ěx2Fb��tl��Y��$ ���^����\�edN\��g�_�u�z9�)���-SbN.�S{���$c�0~��*dY�#�g{��QJ�_�V�o}�q8����kb�x1������B$�֌�O-�:�d�s�]�N�F=c�"���ߟBv�� а�&2*Ǟ�.�Vf�F�ٜ�s;��}2�gӼjk��k����b@\��ν5�6��50��ӑgp�8e[�>�CT0!�W�|���!B�-^��;����,��WR�4}�zNu���4�R�@�Ω��t�����7}iw�:�3m�����O�~�g� ݾ��$��x���@cM�\8fr�J��\]�L|����]�t�#5�"�*�x�N�N����of
��n�r*�����ܱ����3
�XYUB-7�P �N^<]�\-�J�����ͭN�q�Q���� O���db+��)�:�FD�J�1;�-7�=ꢥy��_�jiP��+�r�7��O�����xb�1w�ֲ��
��4,�J� �Щ�:�'V������$h���SuQ��nR�Е!�	���G��/=��(�3�\@�!&�vVOO��=�<Q��ԅZ��A춻����uI�) 2�H���a�LQ<��SɫV�i��v�`��2�?��<����Y���d*e�E�.ʊRW��GY���F�7�M���,���.�Y]UZ6����b��$��;6ou��k��/m׽֍H�1����=d�9�	 W$�^lA���^��6���?�MD�>���\��s�����m��}�,��kp.�z<wl79��� ��;���e��b��p��{�ּmd�ky�-���LfSp�+�%z/Y�%�i�,����=�х�3�dZ��,�~�+��e<<K|5��p�muS��R�.&Ԍ��8�`uzD��u��/���H,:�5=>�">�#��Q�V�Ȉ��~��p� L
���%ub���|��1�+����<���x�>�x��D,U^��L�G�^��^u�P�Օ(j��;��2�0�Xvt<1FS��!�b<��87��&0�ytP��֏�E�W@�Y��Uwf=�O�&Sﲥ�6I�`V�y�z��<�Q`p�е�[I6�M�tr��ڍ]�t[MXU3~�7�8��������Z�˓'��ҿ��l�=/MuyO��EZV����K�|�Tٴh�X=<���R��#�fNjf��o��	<Fr۱E���@g�s��+S�!�'��uC �-�j�R��Hb��=�3�d)�'zlo�"����"���|�T�-�&g�cG&a9�d�C�sl�`�{Տ�0dJ@[gΟ�\��U��[!���X,������N"	u���I/�v$��>? K��9�"5i�~�Nb�y��ʄ�HG����41[jG�/�r�r�~���S%G�4��5��o���D=��9�	1�n �l�����cw���t��B=t����G{��^�/��&��pe���e��)̪H5��v�p��F+(#� ���7<�7�Ȁn4�7��O���*,��Z��+,ӓwG��H�xIy�o�vB�L�tw�w(:E!yzؒ�$��J�J&��g�`�;S>Ձ��P�՗G�]к��vt,cS�$8���L
Q�\ڤ�+5�>���J���F��n�!�v����p'����F鵀�!DO%��?���T��o|��ss�je�.%t�4^'+|��c�ʡ�u�ĸ�w���4��Pʺ���g@@j;l��56� b�o$�=��R��N��P�"8}��������p���4eN<���t�xh���Eg�6�n�2@��rf�ս��4*ʭ��Y��?'8�澘�����:���І &C�:�7uTFdfx�W�J��	���mx�_lL�ޯ�Yo3w���EaK�do�M�j�~Xo��F�F9<.�Z���@�������Xb��%a��A�%-%�{0'������� 8�L!�o�V'�����ۯ�p���<��ʇq���uW�`����N�p�b �=�����6���ո	J*Ѝ�8�QL9!Dz	�t�CF�jm��C6a�p&{1�A���a�	~l��F�#�E�yK+�j�g��ї�K��B4�SF�I�=��b�|P,�{|�T�M�:�3v����,���̓��r���NQ<N�"ɏ��륏\���\�>i���0���2bÍ�x�UP��1�(�;�5���sp��T��|�~r�؊Mi9��?��!hT [RNqJ,��uX�3"E�'H!��C<�p���	BpD��t�x�p-�sGU`esy�&@�x$t�T �����v-٫��ĥ�ς_����{����[�^|��9��s��p9�@�>t��q04s��.�-����1�a�p�̼�09��*/��Ü�5�+*� :	�ݬ�"�FP�\G��[臭Io�˖�߰H.�8~'*Y�4<̺wپ�|�*p'U���]���Qԓ��f�ϴg�U�F][!�(@�'#��C9M�;�'[}a�`�SCH�6��5(̮�"�h��A6�����N��
�C����>n��{�*��=���cR_�q�=��-��	�ͬ_��9�J(����ˏ�"7y�B����/��-��Ԋ�5L�����& �͇kfG� ����Ph�� � �7�la�CAJ������sc�;��b�X_������\L�W���S${m��=�;�,�"��r@�O�m�zNW@��	�v��	Ni�S�����=xE�-���f��z�����GI���O'm-8��ۼ��fgr.����/L؄�6c=?lK�Y&E��Q����S�j�l�;���jp]#�O1҃G�3*��uT+%(D)���ۣ��L�ԭzZ$�
t��J�$��r�뽟�|չg�yO��km0��J���.C)�?��ej%}���w-�>(��z��m-9/+�f}�������f� ϭ͡���K]��[�ca�5x��GT���k���g"�*j$��T��z��?����ci@����>��H�m�u���P��R'����\�]��&P�q�"�@�˲��B{-?Dw_=���`2��\���?�����QŅ��	x(f7sq���<~
���"���;u�'}w�K(�x���a�0�O��*f�I�b���E���:?�v�-��>c���J��w '���D.X��o��oviD�EK��	ܥ���B�����sEC�Of~KA�1a�L�;0K�J�4.KXe�F��bBl��3�������/�c+.:��5��y��@5;�J�%}�B��#!�ݕ��Jފ�C��5�%�Z�&8�������^δ<��:��L���ۿ2A#���|:n�а/�V�5{����}�8�Ϥ��Z���*��f��u+�q�հ��A�c�Ska94����G�b��pl<�����.�ﲫZYQ%��Ŏ¯�ެ�ܤ��Ju�Z�¤�q�خs����T���/�p���{�[�
���E��@s9��5�ek6�ä�5==V6�[
������� �Y��W�Xg;����k��5�M�=ћF֧C9JD��W9D�6�S�٪�C�-�F)VdѦ�ڄ<����k�lJ'X$t8@`1Kf[��^�sa������1�C�������|^H%��}���ֹǌ�~�|q���` �A*�2_ȏE�n2�'dn�&K��̈́bm!�����	�F��ĵE��)&�����;�+\�h���'��^�:� �uU�0�K�~�v��N���6�o��P{֜;<��)x�E�EI����jp��]��#�Y���[��[;�Y���z�۳(B�#�t�6Su�"L�n��\��k�ڜ����_����	QG�r�Rsm����I�>�"���]b����p�⍏�`T0�y�XT�'�a�h
<=�(�
�q�EQ�S�c�6J7��su:
G%?����F���۠�PO�6�\���s'�'��iΉϒnE�S�vOsJY����H�n�
������B�l\����E%���K�婤�iN���J�j��̣� ��擹��p�K�֠�lzR�����<����HR�(�\R���B;���y��Q�L@����+!%G�Ya��ڡg�>��i��c ��3���B��[E��;�T�}3��Vԏ^�ϳ���ݜ#k쫛���v��p��v�9�U��sj!��kNI�y�&���3���ݤ�]�L�T�)�N�uE'��f�6�Ԭ2��
��3�y�b�d+�9�-�)Ri��R�7N��q��}g�=��Z�6����h���$��
�CR�RT2<��|t��J 	Jnk�Ac��l�U;�1�;d#R�$�̦t��� �
�&�[�){݃GN,Rca�'�η�2���g�	{�ة*,�, -{!��1�-�/s�a�7>z��ً�ą�mOD�/��$v��d첷����I�I����`6�o�lb�j ����lC����iѦ4�H�P|��^ڄc�e�C����_m;����v�.��`߽���U˵�����*sB��H3�%�V;x��u�H�R�Eg('!�إx�
0������Q��c��Cae�E,
��DN��^Q��i�s�����	�/�2��y��WG�H'��r1)_�B|'%�ff��,>���v;��v���A'�6K9 x�c	���U�C>�6?~$�r9�|��#���@��I���ؖ�$1�.z���(B1���Z��rnk��J���\��������zܙ
���&Y��20H���'i�m�\�����{v��g�}�H8��|�N?v�+�����,�����q�u��mE���Z�= ��!���^��_�Mxn�=�/�fT�m�/bģ��!5���
�P���P̀�P����]�;�	�tN�,e����E@%"Ӥ�̃q���]dIL��4���p_[C���#��Yzp��ӹ���3�A"���G8�y{�����:+\�S�i��gn�������%����wD(0a�d��c�	¸�V������G��To_�l*���/6�����qR�ݕ 	J	�y��M�Vd���_����P3=*�@,87=>���%*�_u�j݈>�oD�K�xJo�2�S�4H�"T�xrqI�?������YR!����ʜ�1M?ЈO�D�7��]Z)��r�[��I:\A7H�Ș��>2��N���H3�g8���Z����T;�h8�FW�V,ˡ*�I�j�~fރM�8\�B|t|�2\p�(��}ӷ�ћQA�"�e�Ү�\����W�3�E�(4��+�)C5���?ch�������� 59'{�?w���Z<Z_si)��{jCr���0Z+`2t𻽠�e��/ґ���L���J+����;�b�n�r�,� ٤Hr>L��b�z���4<����x�1�G���$e�gF|YxU�	ɖ�,&�.8���__<Q��Rє��Ē��[u�
��v�-�UT�8,4X���[.#e����$9���lV	��/�	p�y�n�8���[�%�v�a�
t�_'9���5��d=N��!BY���1e�f�a����t�:=����N��-7��*�Np�����	�<a<�C������h��;��e��c��nx�Z��T6��i,����,�����b�!Gk�_X�@�w.g��v������rH�r�k��l�'����n �n�`��F�(8�>�΍��dG�e�M�M�{6��3��(39�*�ě%��>���܂d�;���a[>=�����S�~�	F��\����?��L=�g�#�]]����Cu�X�!�{�X�@d�{�����$�^�R�M-����!�Lps'h�07�C����`�'���He16YI?�{�n�,04�Ф���8��hL��1�g(������ye��)��0�Wh<M�ĸן�a���+��&����xCrE>��~AaW� �$��d�բ�E
!�_�8;��F��Xyn�}�(���J���I:���傝gm����P,�)t ʛ��`�Q��.�@b����#F�Lq�����͔�7Ƌ�_J�{���k;���7��z �(��RB/ȡ G��'����U03?୯Pr��(�����4%�7���[�!��f,P��dV�~�+��EA*�X̹��49oE�u��0A�n�OMP�MG?6�B�������.�6��"ڙ�YR���X� �Y��g�D��Ll�w��|��R�u��&yA�-tu�f�l�F�oذ\W�QK֔��U�.5������W'y`z��[�x>ٿ9�o>��0��&h&0�2
/�C[��G�;(-Q ��]����^N3��*
CFƦ��"�Z�b�眑�h���n�l�@�>)%1E���B���AVMZ.��ɫ'����:�-���32&�C������DI���cZ׻��^�WDP�,(@��{B( ~�l4��jTAIN�E��ᾎ���";*u���+�9�$4�Z�ߵ���dI.�!�stܵ���Q��yJg~�z�7���D��$���
+���O(N��iq1��S��8Tt�����G��jzG���"�}�~|�;��Zc�'p���^�`j�P.�jG�	�-���uk�ǽh�4+ɩ���oM��*��'b-��m�%��H4q�U��)Y�U �:F�R��lBk>�N���h[��>;25�����' ��*}������I"��ʑMBϞ��GX��6O��Ϋ�x�0T}�ϥ�ࡹ��j�N2h\�6$���P��� ����Er�vO��}��gH���vA��(�[� ��6B�h� ҉��4#k�_W��E"�w�����w�MX�<d$���Ich����ʚ[o6�O�o�pj;F�s���bx������3�V7/���R�D�m�͛U��|�&>���Xi�����[���Y����C�m�C�oWa�.��)�����[�!��Nq�X�9;.����1����a���F��2������S�D��K#�+ᘖ�IJ����ؕz�aB�W�.�&���ɬ�����wO�$�DT���G����z��� M�$�Wi,�<�0����ـ��t|��ԞP�v��RGL~[�
��Y��m��:����ă2�[{���*��1)&���.4�6�]��U`����+U��ۭ]�q�n<,�Aϩ-;��5�,�5��T�g�u�wLڼ,Ԃ��md�*�w�se��C��h���q/K�=NA׷�u�F�3s~8�{%��"����#�P�C���!����*`�g�]C�ꋧ��G�������Qh�o�3:���$p�b�!3��$;h����|�d����w��SY������nw���5WekXӛI�	�l%'߱[%i*�)�!��e�4�?��4��[�ʽ��/���E�=vϼen|�o�l72ɧNܧ=5p��ˡ��h����.�Z�޸)yY��� ru�A'���]Q�q������j/Y�AU����P)��|���@�v��l�k���
�sv�� v
�-zʆ���w8ĭ�,�������&/�+q�!�<�{�T��0�W���
? ��]2:���G�˭��1�q:��%�V,~�o	�&�:�vce�u��ҝKo��@אV�u���{��a�h��:�s�!�]T��m�z6�|F�ɤU!�+UǾ	=�\+���.^g���V}sdnڞ��469a�d�p���Ϣ�0�����h���e<��F�NW�X1����{K���h�s~pFı�9p�[P���iC+�e�?i�I���d�����Qt��B�DXX܈�#��tZ}������k����?�H��%;Q�W�)�Khf��[�S���WBXwQM�����<heN�lp-?����/��������@ON"`���¸(hB�ڐ0/fU�oJ��ɻ��36�Ϥ�.�� �=�iBCfM�(����7���~�@�0X-��֍=�Y��Lwm ր��+��RD�
z#A�=�kֱX��'ڧ�&y��}�2�\޽�1��qoA��(��eD�g	��_U���y�$��s)�]��[�y��^���Һ���"%)Y�Rՙ���0'z	#��	W� �f�C���o�>"&��cbx�x�S���@�Ե���hZ��}�R���[� ���$��|�|~���ޝ,XtdP
�����c�>�c��ji{]���������k��P��o���!����V�;^ym��PH��jǜ/$�$B-,2Y���Q���{���e���#���o2h�w�~�]�f4ux�*
�F�U�ߐ�� qL�|M��\��{R��'w�[��^s���6!��׬�Q��w�����1ɻ�s�¨}k�(ʑg?(�<�mq���~��Gf��7�|���5h����˹����W�* ��c-N&|�GB����p['�9�����!; '�uO,n�;���!�p���0�JJ?~��fP�r����-��^���"��u���6�m�
q�m�q�O��PC	<�/����5-�d{�d���w4�"-�]�aa�6[��Pp���~O������zԚ�g�2|x���[���kemN�=�\7ıi��s�b��>�y#?���2�ߖg���z�>4!�!aa��[c(���Q�y�K��E{8.��$��2c�PÚ�ue�ٹ�K��K	��߃��&��E����(2�W.T�;�_���~�e�$���4yv�jS!Q�����t�Is�k|-ߓ\�����|�ۻ
t\�.��7���B��%7Thʒ2Uw	���F�-���)74��=V�Y�t��0����(P���7��Xq쇈'�#��0��'�(1�
�V�C
�pNn�E���8Է�)����6�yӅ�5��6�+��z6�˿�"m�3^L���@����������W."��9�\�q-b�;)��{����[5�-�sTF�)KI��X'X}������v�lK�>����:��e�w!m���q��;&��d���<
�7dsD�
܆���,������Yn�1!�����S�\=E����(}�l�L2��~���"�x�S�"/��J*���.��h���,D������� �dD�,��i!��6�n��ӹ�x��΢�<��B��|c�OqӀ(1��VL��6�zٯu����"L��`���Rw>����tf���zZ2�y�3;H�P��uy��<W#aI�{k��~q��#�GA�a8T�����g=����aGKj��q�_���s�zj�U���K�>x��MCa�1m�Y�P�I��[�/�	/S�Ôc�}63i)ǭ���&^�d����ٕ����H��"yά��?��۩?l����Aik+�_��|�4�Q�C���&�����+����T��)CGmn7@�9`�1�T�4~��J+~�GL��>��J�=�A��q��0�*�g��`��G�Kz��n��OÛ!�����0tؐa��Tɕ�4{�H�ʕ�Z.#�x��I�v~����P��� OB����M��rS��>���W����&��e~@%��+ʝf����L�����@�_��u�J@~Do�*�,�5��3�E��V\���,PaY����W�d��5ǧ����U���� �!ZMS�G��5a9 F-Z�B�� DY��a@|�K�Q�i�梴_\v�C�-�ӯm�M7ᖻ�~�Uƒ���3�sl��f�T�O}lb��-h��e�}�R��.�.����bES#����-�y��ƙ�zTΔ�:��6�;�T��3x����V�Mg9ҏ�CG(���e� ,��+��Q;`W��� �m�Q�� Cio���&,}�)��f��o��H]�A���k,(D��֚�<���H�o�����'wJhN|>����p�"�˥p��J�,��3�>w�N0��(�|Xs3�y�"�����E�	�ۤWM����
�f���-+��(Z,r!3�to��5����+�t�k��QsF$��kPeg�yW���N��̠ܺ3�]zxИ��$����{r5����ly��P+	wN��&92I/�~��-�B^W���J˹X��r����,����'���ա��E�2��H~;����U���󋰁x��G�������qi��?#���P��_.�g�}'�O^E�FuX�R���k��Ʒ�K#�C��_}k�*8N����>��о�!xV��ЅO�Z"�������9����ǖ|��Z�<ݢxc���}u���(��č���"�ܑ��i���MH��Y\B�w���̬1��nb�k���C&Lz�x�#�=�1�q�������KT���j�afN^�$���	�4�I"|�ߵ���T�>6�(�灖H-q�b�8Yֈ�-��g� ����;��5�xQT]q����Z�\jLi!&��?��=�(�Ǵ�����hЉ����K o�Bu�?Ϡu����3~�Q,e����K~ۑ_��es� �iU������r���0Z	����n��7�
?�*�o8C�{���N�PY5�/�C�r��$�0sđv��J��LxY9��Ґ����W����-�3�u�`�n?�����S�z�C`��B�ܘ`<��q+$�R�pW�"?�8!뀣VEe~�gn�n�:n:�*Ы�E�T��(�2V:�s�-[�72S��wQ�����I��?�3?�׉��S�� �3ߣ�.�vW�HO�)��an��֌�n�~�t���=�L�҅a
�y�8w[���Q��bѬ3
S���*H�s��r�'	�:k���E�TD8����k�F;�W*@&E}�JFhr2 �le�wY6��ׁA ϔa<5%	�j��>��!��,��20�V���P���%�"�A	.[0��d{k�_xKt��9�=��C:�>�Ե0K�xS�TI�1�y�8?O��$,�{�*c��f��*~+���BAŉ�*�\_�c�0u�RLU�_m�e�)l*��
ܴ��k��Eh��S�������Ǉ�b��i�tȈg����?R᫯Ѽt��>�`gm�����(sټ��3Lu6�'��@L��%zuw%�\�ýne߉��cﲭ	9���� B̵��@�*�~��v?�� ,Tܮ</#���P#L�}����}��~I�p�
E&��H���+A��
0�	�fP��o�EZ�2�s*�<y�PC�A��@�ι��nK�)���es#�Ɣ�_���Q�n�#��9�j]�QIdC'y��8]cS��x�̻p��1�4�M�j�ͩ���`���捽��U�Hj��>ZLj ji�j��R�<D�1�b�j�asZ�';ߙI�ٰ�c�^T Y�������^ʛ��F2��hF��=v��
f�œI��յL�5��k�@�D�w1�/�g�ͣ��o/�ȉ"�<�`�q���~�#Ub�m_\�+)��r��^�^&�R2�Z/B���d�j�� ����3uʀ�c�b�=��%��/�G_4α7�O�o~�:-�〧�W�./�[��j"���zoz8An���OM�(N�X�d�,O�W����L�q 6����8�?}@1@����#L��߁�{&����굨�􌳫���2Y��;�rv/R�0�
hn��Eմ�v��T�Uy���1A���+�
-�a^�j9���
�9�M9�Ȉ��m����ҭpĜx���ȼ�����:�[J
��2A*|c��H�g%�W5��͋f��ለQ�j�Y����
�����S�|b�jK��	R�N��R�:A�|9e.���|���g��[~h���_&!W��Z_
�Vl�a�)eD��Ae/��N�த���b���Y�Y��=O�- C6�-�spC�����,+:bĒ�4�Zi���O�L�^6���n�ۃ�e�6i��ְR��Z���\
>�o?�tcy2�����R8�,�!h�k[y�ɻ4,���^�uꪩEU�t��/%~�Umha��a�n�8e�؏�Tcȋ��>���JIsrm'I�?�Ob7�-w�O���hc����[�����_��a����*�9d88���)��'�v�Ȳ���È��-gp��).�ʗ f������̋p�ҷ�=��*;�9+����X;�B�]jA��\8�hK \�`G�U�����.�1��3�E)���� ����4�e�(45�1&��D�8�3Jo�]�P�'�2���9�]ܨ���L��)[�L��d>rl��jN� B؍=.��]�H�4
�}��:O#��j^ѫM�ѵ�j�!��C�͓7l�#1a.�r� {{�Y�s9�,�+w��O���<&
� ��y~�P��=q�����q-Ճ5z5���y�dyi1��ӕ!�f�#�OeE�T�t�x?S�ד����5��m71���	�d�K��Peч��1�Z�8 �J����f)�e�X�h�)�Q_�nA��ܧ������3)���7i�F�����M@�&��3I��%�_��u5����n��*�w?[;;�Q%	 �&?P:��O�'�~GO�}�V]����^>K~�����u�`����,�0����=�ڤ8�2�)޹���r�9(�	j�?�WD8O$��gR���43����ILo�A��R���c��&+E���h��W�d�j6�������qm\��9�		i@hJކJ���3�Gm�`��>��tZ�<傥�%���иL��U�gj�`��H�oR���5���Y���qld�(����v(�S��^MKB9"�E>1"fp����J����s��8��?Z����{�T ��ib}U��徼z&���I�$kE���"��΁vd6�zm���wk6�s��	Mt�*��'����������z�ֹ�j�XƉ������qS�&�M��LG}��͍�^�I�h)~Л[Ɖ�X��9\ײ`�~}}^�����N�w "����)��EO���$M]�����y�GK�@��o)��|�.��?�W0lD��
�w���O3�Qˍ�ݦ�J��m*Jh2�Y;іLT�'�~\��%�(	 ��WR�Q��.�I7rop�g��T":�f�3n��$�zjI~������g�`3�q���`׊�/b@̀[O3�r!��$I�K� ���2<e�T	_~����-B�P�i�� �ϚX-L(Y��O�r�V�K���^}�%����㯀7��2����~l싧%,#�͹��D����F���T�z�F��X,�ш$����ϝy-
V׹��tO��yeL!����K�����P/#�HIB�rAe2��޴��U�mH�Ei�ꢥ�/�Z#La~e(�#��'F�io�1sQ��$�ΝZ�`���b6��S�hIL)�;��Y�|VD�_s��U{�������~�l�v���:Z���}`�-f�l���9"�o��Ai�Y���l�M��A�qF1$Sp8"�Q���H����K�B�pU�=gL�]s�)Q�]KS����D"�f���J��ԋ��N8�|�|�+NOt��e#~ jTɒ,��/99�w�K�-t!�%&��dK�z��g���"Y�2+T�ҽ{}x����{���M�yrc�H��Jt��%�B� ��:qws��+/�2���*n�n�ؤ6�P��2��5sqʦl�.�e��1*��e��_�n���X���E��6�2�f{��*�$-v��2<d=o�k��4]��@A7Z<u4���ž�vn8�C�rh7�-����+`u��$x�K�Z�vj�m�"#=�m�׫&������E���;����R�����銧�
bxgv�:��N��ܢ��I;�A1�_�tSR�}��d3�YӓޞC�1-��{[���Q���=��-e�x�\^v���l>���
fSX�K�C�ZםW?t�H}3�DzJ[W�}��F0�-P�k�+E�Ȋ�����}�/~&�.H��Ճ�d����Q#�OA�_0l�SwrV���{5w#u��)n��&�`�I\����,�S��1~p�_��J���P�����?m�TI������i�
�f�m1A#���#E��ZV՟5@����M� 0z�"[ծ�IQ�GD,�wxsVz8����E��zQ�O8�,E�M#�Ğ7������H��V��^�����������2:�	e���[O��㰎�`�<����A8Z�,֯joO�\��\��b<��D�㫛�%�ei}�b����8Vκ,�-��3�Be��>uf��:��/�z�:���<���T<�yGF����0's��:ԱlX��P���\3j��p����2f�׀��<]`.�J$bup���fT��4�⛇5��k�-I���� l�����$��鍴')�fُc�꘵�^�����o�rN�U��m�v� �sS�	�
S(+�����{ֆ��hzt7F�Ǹ���ģ��K,/�B�=g�I�Z��LJ�]�_끦�q=f�ץ~��ZHKչ����1����|����8�T������ap�plՎ�%GlNU�4�O:<�n�XU�^p!�ch�;�>�]�'�?����H=�����������Z�odH�:��a�3����
�W�rU�S�2��;{��~_�^r�':W��!��q8���WQ�����X���DM��g���|���Va^�7D�IPG��� �p�{Y����{��̍�x	E�`0���L��C �j���<V8۲~7]����K��V�]��P �bc�=}���Ɓ�{�]�ё�z��aʮ��N�Խ�&0�}91$J����y����'é�Y��P�6�4M.[�5�u9���S�h��+V>s�^m�B�� #��s�������h]�ʤY@OU�;��o��N5���5w�hUo[ʍ�*�}�Ma&ԇSŪg�'쑴�J���f�����C86�J )��GD��Hԡpo�_͸ �,9�&eb�(�*��WVQ�F=@�g۴1��$K����3�|`�}W��|������$w��`��=�4�H�W��8��\���	/R���Mq�»�q)�*��Fi�6gӚ��!D��1�F������P��/5��x�k�f���w��~jI^|�d;/��R�֝5�m13Tkd,�k��� r�S�>s���B!.�uT`����J7��n)�+��.oD��A�<Ato�a,_M���'�Bp�2��)S���Nd@h���$�%���vأ��d`�%`�^�S"�%�UC-KѴ��"~���f�\�N�W����M{*�|����k�@s*��D��s�6�4! :E��`��N�5�����I���0���� c���-�-"�O�19xOXaFh�re-�M=�\2Af�g�[W�>U�?�ro$cbs7/����?"��`+#�����h�1a����̫�
��\$�Dŉ�'m��B��>��FrpYw�=��[3�h5���Oљ�,�ܛU�-�Ԓ���ȫ��A_%$��׷[�X�ƌl.x:,!s�Q��V�w�2����x�8rxG�ٔJs������=�	v7�/a�v?��o����G���� �;����|�(6},b����,�9����ަ$�q�� ��3K�Lm~�w`��(�"��_qîv�>w)��j�����*��X�V�+b�.��z= �>k2��S�3���a����
