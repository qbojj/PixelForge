��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���Dx�hH#��Kv�k�T�t��H ��1FJ�J5 gB2��� jNtVB�Bn9:�M�+Pn���T=�\ɓ�k|ݘ����QV�B�玏�t�R�vz�_F��[~��f�a�;�w.�<z�����O�1F{���a��zh����;�.�atkh��1��a�mC7�����AQ�sw���[h���q�s�_.[̏�ġ�������Y+�PEA׌*Z����@����k<��
j���&Y�6UGټ����-4�n��A/Ѧ�]��VE1�u,*y=V*�0m��>���f9��=��~Jx,k�Xz6O����Dʶ��y�Dnc,g}�`[��e�b���	=J��lY&�YQM�-�v _4�t&P���<-���K�cfq�7�����|��+�9��aQ��� �Y:'�p����Q=���R��A�*����fS�SZb��o�x�3Q�hLg�M�9���D�!��vM�Jj'� Pd�R����������skHN��.j�䚷C�
�.q\_��נp�AW���M������{o�5�Q�,�bD�ՅG�n�3��� �K�t1����
������3��|��E�mp�*�7 ��l��Q���*����-	#���8�TC��`�w��h+�:*|�Q��-�	{���~[*t��=�
�ȸ&a�y�\�j�x��j�BMJx��d.�������%���Wo늩K��x?��3'�ek�>F�)�lO9�� $�#�?߇�u\�A[��
�7g	��i~�# U:�̴Z��z���y�z&;|(o��I7�� �Vs�|�aWk�����nh�D&{�nn�sʱ+���:P(1�DY痷��#׎�]�a_f�ƃ� ��e?Z&�V=~S;���L����"@�"�\���E�C�.��wK�|��'G��z˦0й�����*���-]�xձ��DW����+�|�Ӄ����u�z�N�QAz��U�j���`E���/ B�K]��?��@M��0�޽�2� C2�t�R�B΋�"���l��2Xu�迊}��F������* �ܝ1�p�^OD��E��	Q����ȿ���4NHX~�̂2T?b�q�"{���=K�Ա�Fz�Z݄�w�t�<����JM���4���Yȕ2����b���|3�m�rxl�@��|z)��6!��u ��Q�-�	f�lk��<;\����[H'��Z��h�V2!)>qau��O���R?K�7�c�M��҉��w�l���@��7�]PN3�vƭ�L�ܣ���K���(�6�Ԥ?�*�a߇��q����iD�ߟ `v��RpVV�"�wMS�i��9; ��Q��M1'U -.���.}ha3e�;p 5���9�Yz�����fp��S(FN,�TRТ�=n=.�odԢО 6�����1�5I�N/�j��d�/������rW K�OB�ܫ�˿��{��N3����_i�v'm�ȼ�����T��S�%e�$�o <�)9��n��͡O�8U�����~�0���-Q?�#�����N�k
��n�l�I��Sז�^��=��>��I�zꮆ�YhUͬ.AAs%�/@� L)�?D����k�.br5�ޛrGF|j<S��A����E�r�=d���[|�=����� ;zE�{���1?�ɢز�;�`����G.+��Qq��I�����΄�7ƨph�h��r:�:��M� }�yђ@%+�Mƚ�:031�6]1���8�BHGД��&+�,��E�0�lj	4�k[8��X�y�1�w���ܤyu."rC�=��W�>���0��_�c9#P�]l��E`?�=���[N]؅{�f�q&S���@7)y1"��䦑E�č�^�lcx;8J%g���I��vX�w��C����Sy݋Wp�����.)�E��P�
�,���w�SU�!�'��߂{���-tU�e�gL���C��~����2�^�C}�&���Eˠ��e08�y9D
��&�3����D���4�9���Ai��+{�������ؿ� l��G� �^�6��N���0(�K�Rف>H�Ll��N����n�	k�s�d����x���4�N�y�� �>/�Ƨ[@�\ \��O�2�8�1�uG�%�_�}�э�\���ß�v8���r�n[����Y��2��kD��Z�4g���j<`�(�\hC�Nm�Q2�QT�������<w�h(��a�ރ�+���@ Y)̏C��a�Ņ������~�t_��J�`��̧�uen][s/&L�"9�hك�V� W���ݢ���Z��jE�	��R��9���m�t
�#�8������'c���f����PG����S �>~����Ұ�j�_ �8�?3U׆Q�J�p�t�!o;Kǋ�3�uZ��V}S��.�&;��M �$��^ڱ��
�l4����R8�(L'�j����u��ӂʞU�Ʌ��������,�E;tE�A�\��Pi�a�t_�S�2�3x�ί"{���zg�ྈ�H���l%�aK�Z��3�l�c�u���B�N�)��-ìl�sfetyUp�6�1��gn��
.k��U0�7K&��C�aQ��P̱��G�7bSW�9�&���<i�k��|��ڵ飉��2���\��s^��3b���%D���S!
NM�T���CG$��Q.Wߧ���V-���g�Pg`�㾋�~N����
��k'��FX�Lz���^���}7�K�.<�^!m,Cn<�Ж���vE]�Ԛ�W�U3�"I�R��q����Ò��-���M��TL�4X�k@�(H����0
����np����nT��������v�y�a#��F�cpU��tp��5��
9#�5ޘ����I����`%��|�Ћ�!D�{�X��b���k�/!�:6$)x&���O{�nh��}�\�VoYu�}�)�
���!t��pr�ŝV��a�q{C]��=P�V;'R�,�ݿ�;�.�-��\�b�v���ȵɧ� �ы*pJ�s��e��G�c��kj���Fz]����q���^o��h��ߪ�/���!�����])�V]K~��J�~>��@t�sC ��l6.����%K�NYN�`��]vW7�6���#U5x�?u݊u��ϼxx{0��w�����_��L,(��X;1�>3��?�8[,V�P�����r}/*��g����K��VxT�qqN�i��.�-"�K	��!2��h[���^���PJ��{Znä��ct�)�Ȓt�r
��/��6ɒ��c�n�d���f[L��� <^�-Т��G��v����S�z�vM��s"�\� x��c�	�PU[� ��R葲c���D�
���te&-�x�e_K�tJn�՟�ݴ�z2�5�H6cb�+R��c���U��K�Kr�tp���B����.Bn�ި�����N���p{�6�;���}Y}Z��Q7׭4��W�C{�w6k�ހLO�ol�`��tcSLl�Qv�:H�=��ڻR*�!u��AXh����r�e��.tUX��>��
-����X�зE������+�-w��X�7���E��QO�ht}MG��q�l�a���d�y:������K�U��H{��jO"O�DF���~K囕��?�����i���$����7�����b�P���A��ުj��*A��#r�KX�$����h��<4,�WJya�ܬ����dz���Z4�jt?��-��2�1��o����ǥ�B.�Y�l�\`�&�`����w�T�����>��+bmo2-1�C5E�u_3����?�^,�����Bo3*?Z�Y�������� 5��k��=O�����R�]�j�E`#�!�f��Y�y~oR�g�\M�_��'����7J�Y�xUtE`���\t5x�N�Wˊ?�C�����~��d��`���f�a_��h��>~r���y�lO/���j�z���'F���*h6ۛ��z��ԍn8�}N�w4x��m��;M��oh�ƻ���`�٨�P<��?SI���'�g`'$��3x��R�Q�*w��m�.<3v�H�ʢ�~b$$��w��$�����8Bf'�Χ�Z��x�#��YuR$<��	ɓ����#b칶���Wh�ZER����ߞ����<�C��W���l&����<�"lu��ĵ��Q�cU8��.xCKi|/X,�'��%����F�:3wOiɈ��i��`�c����Ǟ��w]���@"�s��^f�y��F	(����J�IR>d�TC�LH��<�z�sJ�K����A���+�[���L�������b#`�F�/2�p�	������MBGk<Y��f#Q;%`Xֹ5S�8��[F���z
;muy�8����r�.�@=v��^`�4-c
�T-?��d����$F~Dv���p@�����'�f�
�As�QC_ٵV@
4F�5n�k�}��B���o�F[�.V��X��RٵR�������'aO;X=�w�T�k))�8�(��nF]W
����nf������[b�ߘz�`������t�e7 }��1ӳ����0����7���+�]G*��Bj�h(G��+�J����H�>%�~��$!S܇7]�J^n"+��6�K���B������������R�-4��2��찛��������v!�+�z<�P;^>��H;����*>U�t�MU���TB��zA���$�Ba9dG��t�="�m��;���)z��P�e)�¯�(���x�yd�7Xc/�=f�e��C��v��@ъ�Ї���Z��9h2�
��).�f��
�.������ܮVG4��4F{١O��ΨY�B����6qi�������4���RRև[}�@�"����q ���6���q��������q�@T��/xl��Z����Iڄu�?�I5����7Yy���]��zP�����F�rK��~z� ���Ğ�&��	a\��w�B�aM��m럲Lm �^�Q}6��q�żt��c=�Ǔ�e�a���d����(�!�����׬;j�[�#��
�v��~Dm���ShDz]MZؿ#�<�%�L!�/��X�KI�@������RV�{����f�i��1�: ��쩣��l�?!qp�q��b��	Ko��\̮����1����^s9#a�i�e�[H�c��i���\������sX}L���$�{�� �PdRdB�v9Ü�uj%T��}zBz@�N�B/W��M�Ѩ��w�d�����Uu����b��~n�il�w�qBR�z�(4���2w;��ȃna���rC�WZ� 	w>�H6�	&� �:>�4LA?�cwV�r�ٌ�=�������]"P�zw�-�}��
ţ$�$%e�qgR���N�W\�=n���Z@�'U}���8:N' ���ݶf?#����l@�q#B�W����j�OQ��p�����}Oo3ws�7PC�FzS��ʐ(@jjx��nA�ٝgгbʹ�|q�uR>�[�7�i鹬�m��f�*h$����z/��w5��p��#3�� շ)kﺤ�PH��[Ҁ/gk�n���&y��'���	�z�%bp��+��_��eO.�sV�wz�N���i6?I�ɼ���W�=Х���-��u�������Wn��X������t^�zU"mBc%h]�z�ĳI�όu����z�%��ά��n|[`\�������~�k�>3�t��l�VG�P3��e��MY�
e�L��0@�;��q��[]�s$��a�����E�v���np�����0��qV�1�=�b,�"&T�9}� a�$,�d�y�q0�bW<+����d��o>��/�8a '� �I�yC�q��9߬������,�|�+���K��Z��,�F}����m·�8�Mýx-�Q5Z�G����H�m<	�H/Nj�&��r	�|�?�����1��,����	 �d�©ꆕQ�g�	�ߗj9��z������xIT+�{+Y�̭Ȕy��5�^���5[����|��j.���mvw�^�&5[7t�w����\z}��ëhm�K�T��)�>�-�V�^ʄ?u���� �:�$$WJ�QHE����:�T�Јy6ef
��e�?A���5Ibg�Y�����s;7k��=u���{�d�kx�-t�N�\������S{0,��8�3~u`40��p�B2X9�V�7�~��w�λg��ݖ�ĺ�w���
C��W�1a;���*�"W�nP�|4f�����_��N���=���'�)
7��=׺�v��vaB*�f�{!�� -�of=���w�6dr])�M���7J	�{��(B�X�W#�c��-g4o�/�jxg�r=�N;wj1t�o��
���Їz���	��܄�S`T���p_x߾�$�"�5ļ!�HI�O<�W����8/�Ò�3J���$I U��D��1)��UT��3��=�*b&���뀈�r���{��҄������Z7n襍�4>;�*�� �j�hȋ�j_g�ȓL��/�D,��Z&F΁���ș���E)쐊 Z������d�r��n�8�e��Lq���x�9����7AG���S��E�}�SC^J���y��Y���v�8��|/c�s7�-x��a/3���8��	�=jU�#&ƒD�m
�q�/3�p?߱|Yz�R(�e��D�R� ����,���-�xx���j�~#�s$S�����@Nk�ڑo{B�]��������Ɠ�QQ���7O��Y�m������b`��	4צ2 ��M�}L������H�h;��o͵1�K(	� 9��5��'�.p�Y�m�����cBG@�[��sr�	`���e� ;�O3r�G�p�!x�fr2.�<qR)�G9xL�*I[�i��C%R> �A��&3l�5sL�&'��ᷘ8D��R㛴)P�0s~SϠ\�#FUm�����#cY�.6�5�������vC'��|0�iꛉ�v7��
h3�6v�@���ꈩ��_m;(JT|O�TvB#-�R�i�H6mJ�^Xj��"���㬈�;�]���4��ʞ2)d�k�V���s�Ѩ��P��)p���� y&�hU�ȧ�a9���T�b�А��]Vpo�r��昔�C��8ɚ��#H��hW����X��~������s	�0Y�Hgk廙3�q	_ށ|>�/2���f0s���ñ�wA+���q^7�v����80��$�E'y8Lj�۽�33��R-�e�:��J�4MhKf��uwU�&D��p��Zk�pv	A{-�=�H����M��ay
��?[|��2v��i�6u߁�rey������*�z*��X���4b��!,[rs��d��"�r�#�4h,$��A��f#�Y��s(����=^M�	!�1����DQ,B�<��2*����g�R.���^���zbptrR��d�cL%6��B3+_�a�[���v߅�]h�(ԁ���<�Cm02�F�|%d�_Ș�r��5�M����o��y�KJ�WH2F�c���I�IJ��o�Q~�d��"/��Ǩ-�O,��?mj�?ͦx�SZ�)'�%/�p�P���aS=̈� ��m����+jn1NQ��>W���,o�D���l�[�N"��cyV�	<FӶQ�����i���&k�0B Ē��0�a�(���6wj*�B#Կ�wC;�(����-���BE 4(�;��\�F�����%_.l�fP郜�^����O(�n�
'�7�f�_ny�!(��ŏ�!>�D~���r��"4�<w�ڽL=��-�ɴ�I�Q�y�s��feԹ��eY֖D�x��,d�``�����I��j����}/A����.Q������U���ہ���|���ڀ<�Ԝ�r���o�
'1�m�(|��S�A�i�˞�;gc�����T+��QSH�5F1?'.Q�)W(c|�Um�v*Ef���o��>(��4O������>^O�H�1�Z����or}-���o\V�
-��^яfm��E�8g�>����tC��C�p%?�l�Ƽ�����󓿚rv��eB�.1�AO�T�lRܓ'�-@�!|r��"�;���r�̵���6[����tХtcVq���J*zզ�=Ӏ�k��"�V<QPb�)ԧ�{ ȡ:
��J��X�N~�{H�0lg0�{�BN�Zc���A��� �X$�$�)n7q��$��U�PR�e�\�K7FI��~Z�f}�s��F���������"Z�i��kT�َ_��BN5�+I+0�k�\D ��@0�i0b�rm�k��2\@5�����.�������>K��笟Nͷ),|/��o�b�֙@�!��� �g�LR[;��f��^��n�p���n�V�A7D"*����F�`S�&p�}�B��Uˀ�����d��M= �%�(����2��5h(�5V?��������3��eB��1��)P]G6�z���3�k*����-��q�̧R~�qk���/&ѣ�A��픡>�v�0�\���C�2�F����2!���=c�i�ǭc�4a(�b�!�#�����8���j�w ���>�=�OaW�C��	��ʙlif�c������H�~�_��<L-��;vNC��~!8�07~�^���Y��h�����1���l�W����-73���<�,����ni�O�����
�<��2ǼsAϯJApB\�ڒ/\�)"3�]�mc��{}8Ȋ_O$� eX��Kn�$N��	�Qafp4�&^b,�㪓fX�pI�������X�K�nӔ�fh�-7���-e���6�ś����F�J��c�dG��]�5bI��y�3��e�R�mn�_��nٙs�R?DO�̺ �_�!$�kGO?�+j����$�iZ;$�m��G��7̓�D�;n��SC�1�x�k��K޳r/sS�w#bE[V���H[7���E��0��� �4zo{���T3�'J����S�)R��cض����.{*'j9e3��H�T���|��w!Pz��E;�w���	cd��W���\.����_|���kat�t�U�vq@ɜ��%я��'٭��	��BjK���I}`�����v.9U$�@�݁Od�B-o- ̀[|��4���+;Ԅ�N3g�Y*��:����R.��ݢ�^`�!ር��3��3��"'�8h�sË1��x�3��đ���f��w(؍8�j���
�l���f쿰:"{��A��A]$��<�/xj�a�cȲ�s��YiY�u]|c�~��h�x<޿py4�i�����A��$)�bz�4!�S?-?�ٷ*�ue:�гOy����A��i�ȍd�"�R�l���˘i)����J8
�Sm#씦b��O=�����O�}��~8��~��[��#��J���.2b�U_)��j�JK��x�ym�]>KIj�$�`Jm��ݲny������>o�X�3dHŕ��`��z�(�{�NYyҊ%�|��M�aU����dX�>�3���ʵw��o<��4��	�6d���k���"�*�̫��/𕄽�2�%I�5\�SѸxi64�mUܯ�!e�����2�RQ�b✱$��e��>�/��6���q���&d��r ���.C�����9'};Nӄ�����4�r,��G�zF��Ae�;�od���������܇ݔ�6�W8o�u�ت�B��΁x�	�d���4����1>��3"6z�����`Y��.�#q�i��}m��+�u	sG�b!�m�-1�ȍ�Pg�E%�u&����8���d����$q��BR��-��&|\4#v�֚9���(�-�3g_[oS(g���zrf�j0��N0l_���1��9R$u�Kw	v�v�@'0Q�4h��X�3�����Y,�����d���G��@�/c�x�?��ch�?Ȝ
`�-if���5p!~�����Q]RMb��̛���!b �V���q��3
�b&�[�M/F�׳��کw��)P�����k����?9鑝�I�䣸%�h+���pG��Ó��4O�nyAӿ�{�r�.�}I�4|h��:y/��~s�^8��X�r�� �M�}&�ǬѾ�p*9�*����/�8�O��M@o��\BoQx���U�3p��9:�v��:@x���T_Dt����~�-%������F^2�-����h'�K�����#O�?_AX�
;��XZ�Rh��T$�֭돜��(�bA}g��5��8����w��i�ÿU�m�~�QHK �#f��/%̶M;j��s�l:�6��t���!��=>��&�/��K�Y�QFb�{�7��x���ǌ�O�Z�ZU��;��"mEm�<�)�A��&H5�$n'z���و��j��?�}0��!Ԝi�X'v�v�g��jd �����Ĩ�]t��3���
��ج����5bc��1��X'�~�M�n}�©VE��ko4���T�G�4�K��xБ�-��%B�{e�U�i���qgyD�H>� �M�>a�2��������ט�o��m��+Iov
���*�vCĲ̮NH�e��b�fjp��S܌ۀ���p��ّo4L��c�@δ���;꧋�Z����V�˺s<�%���c�`��J��߫+Ay��R����&�f�h��r��ϏE�d���Lo��O��(�����ct�f�����/��¤
�v�Qߦ����C)��h8Kf�'�\&�f�O��\;�����K�s�ɧq��#K*�1zn����,�pk�<���O~qf �e����L���!➏�޽)L���:6)����/�D���hF����Mt���i�S|h�r�ml{��f�]9�7'ǩ��HP��>;=���9y�~y��ƭ$�K������w:f�_!17#���cmb�Q�+6?QŮYu ���)jiH��q�Rt�¯��n�'(}&ܱ���a�
�Z��Of�\%����3����´�����d�Sv�R!�7�!^D�/��/��O� F�!�Ș�p�]F���VzW�Ѧ�j�2d�U�](�3��A�a��jK9��SB�6�(�s:��a<��V��)�0�����mU�R�(Xa������W�4.�I5/0q�y��7�[~�m\�?��,��V�BӲb�#�h���*�ymk`�5e��D�ޯ��>�p6Q���pR�%9���Xo��f��'?G7��m�����~��Ⲝ�sd�������I��ؒ�׍rL�s�"ú-$�
��)��7<�����՝�O#���O�+��)KAY�����B;`ޡ��ˤ�`!5c2����D������@B�B��O*Z�k�E7ZC�	AݐR�$�؃n�R�)`P���Hn.'���-͛�|�Pd�td��4YW�Z�K�#��W���jSz�����*n����`�*�r_��:p�%X�_�+�ޞ�R��u�l����^��1��
�SeB�x��y��G�s�%PP��+�b��SԾ:��3k>iI���Co��.dl�eTl�A-�fe�`�ړ���k�P�ڦ��y��4BOx,�UP�(un �P2��*+�G)���?b�E"�-e6��������7�4P�/u�mL��5)�݅b��ԩ_9�˰�=o�v�)�m'F'� F�!ԭk��m��#����i�����5�G�������a��|�=����C���<Y7<(6ƳI��@THz:Q��F�z�1�xV��y-s�
�A�(8<OHu M��"Y ���·�N��q���*X�sN��N��\ct�r1��ka��+�I0Qf�
�$� �@�".�4�4e�^vmE{+�PC]�c�����3�۝%���&o1#Ȣ��n�����Z^��HE� #����ʑK8�o�ȣjd����E=-�����l4����vsd޽:d�}H�i܇e)(G��i�}�낤_1�$?h���g���l��:��̭��qP��)����[��|~-��/e4�*k��Wr������`����r)OYi�����/��`9$Ƀv)J�ZOBF{�8�/��^��	V����+p�_���\8ڎ�{LK�����1�80jᨇ��V��Bq�(�I"���A[�Vx�R�F`ړ�Z0�Y�� ?�e
Jh���E�T�NcW>�ف�!d>�1!�A�:</����#��L��Q��4b���L��I�MG����W'�j��BdU���Ξ������b`����V���!pP�x��?B��'���)>q�;x���e	c0][�!�Ij�i�rG�c��Ί3t�81-�Ѩr�\�f�E0���,�k��ġd�<>I)���wcD�d��hꨝ�N_z`��r�A͠*�K^��q�.���*�]�+��̜�yU�'ZȘ�D!�6UK��fc	�p���+j��Q=���i��J1*�^�t[�PDs�8�9�;g�.B�.�9�q��l:TL])���^��T��h����cp��iT�:e� �1����	?1��A��8�b��(����:��p�������:`SX�X���Z���Z~>��Vy�>c"�+�i�o�l���U�����$���2 o�����nRa�;b���� M��Us��}�Jr<��/�6��S��(�=�
�3���x̟9_�����E־(E�h����ֽ3���B���\���"�	��K��D}���� ���/h�۔�8+���z6� ��Qc�X�{N��5�K�ص�����q2���Ę�_���p�-6_E�.8�Z�u>f��������+'���h�d��(�G�[��)��S���Q�a3�lb]~�Z@o�ZطJ�5����K�����h���������'�8��4O��~�D�t�l�ހ	1N����R����o�^8CѴ�w<���Np�cy��ҝ{�U0.C�d��R��T<�|��9���}�/U
�C5w9���[&B�L�ڿQ�x4���ẃ>�5�m@���LU͔�
