// soc_system_vga.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module soc_system_vga (
		input  wire        clk_clk,                //           clk.clk
		input  wire [1:0]  dma_csr_address,        //       dma_csr.address
		input  wire [3:0]  dma_csr_byteenable,     //              .byteenable
		input  wire        dma_csr_read,           //              .read
		input  wire        dma_csr_write,          //              .write
		input  wire [31:0] dma_csr_writedata,      //              .writedata
		output wire [31:0] dma_csr_readdata,       //              .readdata
		input  wire        master_readdatavalid,   //        master.readdatavalid
		input  wire        master_waitrequest,     //              .waitrequest
		output wire [31:0] master_address,         //              .address
		output wire        master_lock,            //              .lock
		output wire        master_read,            //              .read
		input  wire [31:0] master_readdata,        //              .readdata
		input  wire        resampler_csr_read,     // resampler_csr.read
		output wire [31:0] resampler_csr_readdata, //              .readdata
		input  wire        reset_reset_n,          //         reset.reset_n
		output wire        vga_CLK,                //           vga.CLK
		output wire        vga_HS,                 //              .HS
		output wire        vga_VS,                 //              .VS
		output wire        vga_BLANK,              //              .BLANK
		output wire        vga_SYNC,               //              .SYNC
		output wire [7:0]  vga_R,                  //              .R
		output wire [7:0]  vga_G,                  //              .G
		output wire [7:0]  vga_B                   //              .B
	);

	wire         fifo_avalon_dc_buffer_source_valid;                 // fifo:stream_out_valid -> controller:valid
	wire  [29:0] fifo_avalon_dc_buffer_source_data;                  // fifo:stream_out_data -> controller:data
	wire         fifo_avalon_dc_buffer_source_ready;                 // controller:ready -> fifo:stream_out_ready
	wire         fifo_avalon_dc_buffer_source_startofpacket;         // fifo:stream_out_startofpacket -> controller:startofpacket
	wire         fifo_avalon_dc_buffer_source_endofpacket;           // fifo:stream_out_endofpacket -> controller:endofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_valid;         // pixel_buffer_dma:stream_valid -> resampler:stream_in_valid
	wire  [23:0] pixel_buffer_dma_avalon_pixel_source_data;          // pixel_buffer_dma:stream_data -> resampler:stream_in_data
	wire         pixel_buffer_dma_avalon_pixel_source_ready;         // resampler:stream_in_ready -> pixel_buffer_dma:stream_ready
	wire         pixel_buffer_dma_avalon_pixel_source_startofpacket; // pixel_buffer_dma:stream_startofpacket -> resampler:stream_in_startofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_endofpacket;   // pixel_buffer_dma:stream_endofpacket -> resampler:stream_in_endofpacket
	wire         resampler_avalon_rgb_source_valid;                  // resampler:stream_out_valid -> fifo:stream_in_valid
	wire  [29:0] resampler_avalon_rgb_source_data;                   // resampler:stream_out_data -> fifo:stream_in_data
	wire         resampler_avalon_rgb_source_ready;                  // fifo:stream_in_ready -> resampler:stream_out_ready
	wire         resampler_avalon_rgb_source_startofpacket;          // resampler:stream_out_startofpacket -> fifo:stream_in_startofpacket
	wire         resampler_avalon_rgb_source_endofpacket;            // resampler:stream_out_endofpacket -> fifo:stream_in_endofpacket
	wire         pll_vga_clk_clk;                                    // pll:vga_clk_clk -> [controller:clk, fifo:clk_stream_out, rst_controller:clk]
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [controller:reset, fifo:reset_stream_out]
	wire         pll_reset_source_reset;                             // pll:reset_source_reset -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                 // rst_controller_001:reset_out -> [fifo:reset_stream_in, pixel_buffer_dma:reset, resampler:reset]

	soc_system_vga_controller controller (
		.clk           (pll_vga_clk_clk),                            //                clk.clk
		.reset         (rst_controller_reset_out_reset),             //              reset.reset
		.data          (fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                    // external_interface.export
		.VGA_HS        (vga_HS),                                     //                   .export
		.VGA_VS        (vga_VS),                                     //                   .export
		.VGA_BLANK     (vga_BLANK),                                  //                   .export
		.VGA_SYNC      (vga_SYNC),                                   //                   .export
		.VGA_R         (vga_R),                                      //                   .export
		.VGA_G         (vga_G),                                      //                   .export
		.VGA_B         (vga_B)                                       //                   .export
	);

	soc_system_vga_fifo fifo (
		.clk_stream_in            (clk_clk),                                    //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),         //         reset_stream_in.reset
		.clk_stream_out           (pll_vga_clk_clk),                            //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_reset_out_reset),             //        reset_stream_out.reset
		.stream_in_ready          (resampler_avalon_rgb_source_ready),          //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (resampler_avalon_rgb_source_startofpacket),  //                        .startofpacket
		.stream_in_endofpacket    (resampler_avalon_rgb_source_endofpacket),    //                        .endofpacket
		.stream_in_valid          (resampler_avalon_rgb_source_valid),          //                        .valid
		.stream_in_data           (resampler_avalon_rgb_source_data),           //                        .data
		.stream_out_ready         (fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	soc_system_vga_pixel_buffer_dma pixel_buffer_dma (
		.clk                  (clk_clk),                                            //                     clk.clk
		.reset                (rst_controller_001_reset_out_reset),                 //                   reset.reset
		.master_readdatavalid (master_readdatavalid),                               // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (master_waitrequest),                                 //                        .waitrequest
		.master_address       (master_address),                                     //                        .address
		.master_arbiterlock   (master_lock),                                        //                        .lock
		.master_read          (master_read),                                        //                        .read
		.master_readdata      (master_readdata),                                    //                        .readdata
		.slave_address        (dma_csr_address),                                    //    avalon_control_slave.address
		.slave_byteenable     (dma_csr_byteenable),                                 //                        .byteenable
		.slave_read           (dma_csr_read),                                       //                        .read
		.slave_write          (dma_csr_write),                                      //                        .write
		.slave_writedata      (dma_csr_writedata),                                  //                        .writedata
		.slave_readdata       (dma_csr_readdata),                                   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket), //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),         //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)           //                        .data
	);

	soc_system_vga_pll pll (
		.ref_clk_clk        (clk_clk),                //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),         //    ref_reset.reset
		.vga_clk_clk        (pll_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (pll_reset_source_reset)  // reset_source.reset
	);

	soc_system_vga_resampler resampler (
		.clk                      (clk_clk),                                            //               clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                 //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),          //                  .data
		.slave_read               (resampler_csr_read),                                 //  avalon_rgb_slave.read
		.slave_readdata           (resampler_csr_readdata),                             //                  .readdata
		.stream_out_ready         (resampler_avalon_rgb_source_ready),                  // avalon_rgb_source.ready
		.stream_out_startofpacket (resampler_avalon_rgb_source_startofpacket),          //                  .startofpacket
		.stream_out_endofpacket   (resampler_avalon_rgb_source_endofpacket),            //                  .endofpacket
		.stream_out_valid         (resampler_avalon_rgb_source_valid),                  //                  .valid
		.stream_out_data          (resampler_avalon_rgb_source_data)                    //                  .data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (pll_reset_source_reset),         // reset_in0.reset
		.clk            (pll_vga_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
