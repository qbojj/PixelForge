��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��sa^s����Hw�9�k, d8y�Cl��7U3÷���@�sZq�W�<*�K��J��h�mS,G�Vs�VM�t�w�������U���Njـa<�\�h|��&7slZ��w><eK�.(��H��x��$<b�3g=�f��x����:�V4m��AWpX}m���&�(�bTb���%YW��T����q��ig����ad}�9�N��%zpg�-�l�N`�T�5��ak7[�gW8�χ���n}ኧXw��B��"��.�!Ҍ�aL��$�Z��2�[GkA|�+�L*ˮ1���U���H��G����Q)N����m̀��0�F���*?}����'KP
�7e�]:��L�,E�k�I
S-�񾘤�W��$ ��f�&f>�D˴Tݠ�$����a��w�LYTn�|���� m|�>�v/<@Eܵ%�N��Ih��r>/���߁�����3C;��������s�������3��Y�pg�|K|O����D!L������o�D@��T|�ǅ���l�/�,��cQ���^V�o��l�$d�y�����=��o�28@F������.�"l�~=�a�R6���������ٵ`�h��u��]�ر�2ScH�y5��ȯ8{딄k7�7V���CI��ab;�0N��=V?O�"`I����ςi��d�@Q�q��@)���	}P�\�r�_u�Eh��j/���;Э����O��	�����H�rHJuQ��h�A��(N$�3��J�RN/s瘬���!����a�3y�A
�aNv��/�載X0�{�~S蕑����9�s̚����7I�Ӣq1P��@/�(%M~�<P}�]SuE�@��� yq��u�7]Cl�UW�>�R�V�T�35̆d[�(�9�w5��M�Y���R[��ه�Y+pw��b���*tmi���UI�&`�c�ӈcɿ�ܸ�	V�~�LC�\F��GQ���2Z1'�Ƿi��b�O!��2i�H��፧'F��-��@*�����?+�?��/�̓�7F]�U/�kG1'H*��Z�9 �٪U�ڒNB��Ǭ�g>?������_�z����B@�'g��"Pl�:z��dO@��ty�3y�"u�ys����A3�ۃ//@ܳ�s ����Ӎ�H8�Z��hv@-��=>�x�b��.�F�U+&���>���|a+��8'%նj��x��j-:���E��NeE���W�h>+��tc�;�*�_��_�!q�)����4Ŧ��8:XTG� 3 ���)9�]�Ia�1g�M��^Ǖ8D�5�
̾��F�����R��L�����2|x�Z��u	4���AdM02&�]�-������V�����D�s��e![@��XI	�:�������1k� �_�0�E�T��0c߭Dkd��*�w%�S�w���IHX���M�8�Ψ؁'	mVi��Y�ni�+R��m�P��ָ@W�O"/�3�:Q�G��k���CFL��9+"��D��4Ak�o�lA��g���O���LWtO�hv%�`��_<��oA��*%�z�|�[��`3p6i��xESj<�(�N�3�ϟ�A*�N��<*[��Y����+IJ��;�3
Yj�+ۤ@PE�$Bd��R&Y˘�Gi+�Ͻ�i:PH$Nـ����B&L���Vz��@����p���ik�\�&��x�A�׵�����x��僾���5�*�kJǭ\b�X9�_�ŝ�(>�a��`�m�3u�f��f�#����5>�W�/,+���`�C'Ud�yPNߝ|C'=��P�,�-w���۪�0��j?��}��������O�Aw��h4�3���8K��	�Ӫ��}�����3��3���WwIlP��O�-�$���|P�!�9��1�ŽoC{ ���� 5��N�.�r��?�A1!�g���z��;0��zfhg�F}��Z��߀�jb�~l��C����4�l���e�Њ���x�������- �q�m�����K�����ɝ[����T3ms��N�lj����<�,g����0\����H+���k����-AOy�q��
T���9�ӑ%�?����/�*EI�k�rw��t�C��S1x�4\�-��g�Cqiܘf �z3�I�%"���|�x��<4��ʪ���4�S��i<^�!3?�w�K�g����v}�ppQG�l[t�?-���"+--8�h��g0ec`��%��+�u�@}xYȞ�c��J����Aj�r`)܁���P�����F\��u\P�+�A�
�g]���+��l�@��UB)�W�FKZ�P�s�W=l�c�D�J]���[��|p�7��fTP��4`st�L���Q�1V�(�|Ew3�6�U���(/I�����7�e��/�:1�3��^V�G�W��CpJ�qx�+ֆ��v�N�|�ȿ$��0��+����{���e3[�M��7(,�f�A� �c\>=�"1S�Mt;���x�'3n0^���<S[�mo��[���<����z�:�WR �u�D9���B�i��B�,�HX�%��^ק��|�a�9��U�S�b�8͂%0rcdTG��>$�+9��=k�\/�t�p�ƈ�?����Ħ^�*�#����Hj�J�0�g�1}rWy�<�A�F7dɈ��eq+xPͥ�S��vX_ʎ"��H�ٍJ�=�;�����F�������K�!��גS�'�g`K>5S�ߎ [x���]h\l����+T
u_����RW.~��:Pk��W�7�~
Tw��A�#4%���1F�H��k��]ϵA�^��K�����uݨ^�Omc��9>{�Cf���0�gÞyAiFW�a| ��&`89����;*Ƿx9+�� �~�͋+�)�:��so�諪O_A��a��,�w��	n��d�uS� A:�Zi��z��?;�Z���y�w�V�e\�خ�G#��d��9�-}�����gёtj���>�ZP�ޭ�i��]5A-?�ꏫy�TS��URP����x�92��F�����=�S�k��m���	O9l%]���n)��Z�7&�u�_H�Y��瞽�7.���#���1�c�� �� �L�輢�	3�sv�?2��T˿���=A� >�9�����_�`4sG��1&/�1��'�
�����7�K����"yU[��:��9t�v�R�p�!���'1ʹ?F��8�=����x�tdv���m% nI�h�<ݥ��Nv�j�H�ˬ21��qQ���һ",�Z'���ظ+�&����ڍ�M�����s��v����a�����������b������ɚ^)@�o~��Y/���hg�vowÑ�_��x{�U��#��Ղ� aXoAv�hݽg�F}(X$��^�j�|H("c�v�-P��
��J��Nd��J{<��y��<�/H_���hO2�dde���Q�FOE���dn�e��Dţᇐ��f�����W�=�8A=7	N���P]��%�}"ӻ�����aT���v3�����|ǅ�Z��cVTf�Y��ޓ���ʂk���������8�.p[%��L<��1�x6��"���9�e�t��;�5j=mdXx�$P{A��YƐ�[b�D���6�y$�c[����g�:��oP�"���z��IT��?{x���m��D=:v7�!؞�7�o6[��yRn�Z�p�5X��ءZ���DP�m��߲�MZ4�h�`��������\�M�X�%3��L7FR������|�a�.�[����r���[=��$'2/���Q���Bzw���h'�ؠ(y�&=ҋ��`�KY�IL ���ɖ�YKr����j�Y��t�]JP�ʌ�p>��o��,8Y��w�9�"�,�ڃIzG�ff�5���5��j$��t~�k�b�}�ڙ������2�J�)���T�g��9���0���J<-�!��>'b3w���
&?<1��%7���֜ď@�㲊�@�Zj.���ٰa�3�7O����O�g�X�	C�,[O�u���y�ƾ�#x���l�Y�@��g����H�{�%,f��ITCw�Q?�zU�nx4G���N�.]$.$(�:�����]��U�7�j��ۦ��_��*y׭�צ�Q\�#Q��m!S�\���Y���]_C�?���/�i�}�פD�5��]kt�m�.i]��3�y���_�;�A�|�����g�bi�.���\>�S� g�:��`�̐M��І���܃l,T�����I���o/�M�� L^����j��u�"n�.��P儾6��/~�WU�Z{b�L��'X��+Iےݒ��VH��=��bz�CNS�m�LI/���Y���.:�����ũ�1-?��DP�!�"u�eÏ���S%���8��>�z���[�����:8"Z�zY��'u<���UW��	�9���an�6�	��q�s�>vtȟ�&�*�g���wU<�4x�tʸ�i��3;]"�U���w�d`K'���SG��$@z"����Y��iऔ�`y����5�9M�1�}82Y��$�Z0a.�nu�}��y�P4uf���N�ѹ��� �M�P�kv��|q�����S����7�1w�I"g)��b��'+�I��K�2�T�8%M�*N��m��X�
�\%�FC��_ �	��\�X����e�e$LRYl�m�x�<�X����k7����tk�S�#�*/���Y���rF�r+�}���>U+�������PY�^r��p���Ge-U��Hv� ������<D�ō��\^=��w���* xg1���m��v.����?���r)AЖ�^��uf�*�����H=���E[�ؗ�ɞ{.lF���`��k��c��Ȕ��E��4�S|��,{�r��yZ� k`�;�p7���n����ґ�۳�ZSԀ�߾�Z���W�����Pڹu�f˶t����Z�HY������AӁE���%z���!4l&�ɢ1p���ծA፵�<��	���2�LW�m����]K91�ּ�T��(V����R�����:si,ӱk�p�poM����C!�HTN�!煟�b�v*>�ص��p��H�PRu_ae=�-��.����糂M���~��gc8��3�]a[V`��
�>��C���{�3��-��l��CQ�1� ��[��+�sF0�ʁ�?cp~\������vô2���w�ek�n�߽�Λ��r3F#��+`�]�aٲ�p��h�wЇ����;<�z͒�����]H@��b=�t���$r$B!�֕Q$L��CV��Hn�_�eǑ_i-�\�+홓5�ɩB_i�G�Z�6
�𝋦td�"�U:����x�fQ��2m�r@8L����R�)��~��8���!u��)sS�#�ϫ�QE�5Da���<��\ҋÀf�T�N�m��W� ~�i�"��C�Ê�1�jI����j�h@����,�B��lnr�Gd�]o�>� 8q��|**�pB�C��;�u��urbL+E^՚
{�P����̎(��#Ӆ�3�Dz]�9��JL@J~��9���b�ڛ�z)�@2�/�)�2������<���*�8Vld>��c<w�I����M+�	����m"��\1�i��J�by�Ǟ���y�Q�)����Z��<�ɲ��5�����xe=���y�ܟZ�������%9�3򣾳��A����	&/�(�j�?.�E(	ل��p�b]�j,K5.{�57���,@����Ï�Q��:W \�S2�u���p����I�d�#"��Xl�u��c&�'�B�Z�MAb�s����9��J���Cg
݅���hY��N�e>�~��x�|N��Di;�W���%�N��Ř �&Ö"��pp��Ƃԣ.k�q�����zv9�I����Է��7?���ϫ{�Sr�:���k�)��o�(B��REД�,!&�`^ԤK���3�!?�x�	Xχ�$a�_nXV��5jtƮ;���P:n&�p*_�9��CO�8��d��@'�%��� p2�t���M.M_�H 0@��-���:�tZ[���9>�\�i�a�Pq�R������D�d�}eB���z�D�Q��@B��']��<n�ӖE	��F�&u��g $�ݖ�U��Kjȩ�D6��2q>	Z|ʧa�1]���.e�{T����dFP�T&C��
U��>�p�^M��m�K8��]bb~Y�=@��>��������n��,I܍o���E�3z۶�l�;/m���ږ�8�����/%�oJ��4�(b����j������X�����돶�6�U�h
�U�h��
�:���E)�-A����d���`�T�P�7�����������L��>�R�U���c��\���l��H�bJ;T���uu�l5O��|��r����ac)MG��W�\1��lt�T�}�!���d�o��}���2�	`�aM��P���J�y���ZDi�ȱO4#�^N�Ɲ���L�mO-�]��U�	'�P�P�lU�X\��&��Ƀ�p�%����~���ǽ0����<:>,I�%�k'�rK@��
�j��s�-U	�'!&7��5��* ���c��i1tC�����~�%�~dg��2�^w�G�PZ�^<1F�.>��,ٌB�T��u?��4���v� ��#�g�)��OJ=�	��G��M�&q���r�՞�8��JV���TV�d����_(�1�9F��2��z�$u�Y�}���G���T�3)i�qQ�_�`0l��>�����J��!����Y
)���_@�;�D�ڙk����V���c�j����0�QxE�f��M��:3���1?.�� 4Uک+�����y�`f�ޝ_��m�y�2���߼טΣ:��?�����FWr��R���Ð����n��w}c�k��]DY���3J��*�)��7~�(�iȗi8X��|��%@O�͎b�ki���w_�:��ڨ9��G��@�S��|��%'}8�w� S���i̒��*���ާw����hE�/���C���6Զ�ᡚ��}{`~9��Q��|����J��т���R4������^L(v }�������~�����5>��gK0��.��C�S��.�L[��5X�&�E`�A���i�e�	ʮ���=��(��J@%�*�uԩ��0D9bPT�����h>�2VX�^�����kS^���G�&Y�F�ۈJ��z
���\�K�_C�[8�DZ֝�Eqj��
s��u���gy��P��`��>X)n>A	��|�f\[jɱ�r�Z��&����e��z�X��&~���b�����/&@5,�T���t(��B�+ZDz�6�M��?�<ʃ)�xA��Y��Qw��Тq��3�|y�GInRE��,ԍ�'M���\���\D�2���T����	�B�/ϐ ���Y�&�9p��6:��G�$�I���"3�W�s+h`��(���3�O�_ɨ�׏΃���+E��+	ã�Aݏ��hL�c�w�[���EKk�d�V�ә�U������=�����F�����U�+ӑ�7<ګ`c�Ɣ� ���L��m�o-�����O2#�.F�:������<�����[��[��qR��
o�F[�/彇��E��d.�V�����SV�ʕZ�+�4�,t/0����M��%��"i.��|I7�dH�.�_�<G�ID���v��{јEz�E���⁗��qڪ�W(y$��{�P���x�/l���r;�b2�<@��I�Y-x��o� +�7�ڼ���Z����Jj���9��D�ξ�5|yQ!~Wp���Ne��xM�o�N�OL9�����	Y⚄>�M܍��Ĝf��iy��t.�Úzت�e�^2�25�~�3�dKA���{�Ss#�Q���e;��8R�Ə���Ex�N��^����V�:|���Q��a��5�ܮ6�54`��l����1�D�[�����t�!�Q|�ֈOʙ)�d:=��8s.���5Zi]V���Y&B/� x�|x��Ǿ��_��ƕR��d_��s�k}�<���mWrPi�P�xu�����Px��� eQ=8Ů=��T�b�b�/�4gq?xj>Qo#��8��lDy���p��t�����w,LBI�I���t4��w��&ݳ���C�1+���X����5hE��5U2g}9����b�l$�?(��K��mR٩7M>�9�)D�.g]�n���f�c�p!��~�d4�;_�/ƚ[�4�A%ޥ\�f�cK��[ܦ�|"�d2�n.�I�-��FO~H�,ӌg�sԘ�,]��=���|�R��
�πI?I���hI;�n����ū��"�7}�;q���{Ga��ov]w-��p���"��!���g:f�/ ,�:�����ۆ���c��/���.'�05�6%��P����Y��,Q��V�N�oۅ��������_i3o�o0�s�;#��|���,�(]i2�vd��-D��_&;7�R�g�
۲P��b�x������AH�W�ٺ�vq�^����=��ӥK2��!5�g5���X<2n�B�v@�EбP�Øm���ǀĩ�*��#8ݟ��M(z���wy�u����?W��LG�Cv2F�<Cbe?Wo�ItWQ]�>�ϝ��CGꞟ-��b�|qn��Ԭ	-��I��y|w�kMh����[��i�D20��[8L�[NИ.�Q��Z~��8���Y��;20�yG����²T�`k��5ʊ��g�H�]�n1��Uo-b�����GE�lUJ�$�|����>��Oک�el8�r)�E��A�F�(i�H4��}�������I��p�?k����S
�^��G�_У.��Ɂ
S��t��t��V��x���%�O��>V�5��
�\��W��Hò��kLʖ�'�zj.��Ӿ�ᬠϺ%�a�[z.ؾ�^җ�qç-L��@�=�BL8C��7���l��Jߢ�g��.�1١3%��3�Q7���t)%�վ%�-�gl��ܫ��.׵s�A2�:��Jýh�Fb,7P[^��o�tԬ�=�f���8fOK�1 �Z��'
�r$3�Ae�������P���_�1^h���_��?zm�O�-Iu��{ɀ�y��l���8�)��<,gr9J{�D�8�$|��pAyČF7D^��Qb�dz҂m2�j֢�	[��m�W(3��N\-���sR�f	���XH�ϙ�U��<���V�w`�zS둘��ɯ���A�%0�,;@��d�2�o�U'�7bT�]�����{0���wg0"Bfwu#o���VR��R)�E2�)���B!��mm�Y�ç�꾁��9bG��g�ǔI�4Ҙ3P�̗�-D�- �pa����c%�5����+8��Lf�ɍ��GW�����hgfZ�N*��N�2p��S�ʾ�kL i~(��4�ఆ ��&-s4��ו⦷D�cMQ����K�mjp�$��;��d�"Ԩ�tf��o|�9{M׍�/�	C[꾲�J���Uvr�/�	���FlTΉC~Z�f�N1������K��HQ���.;�GW�6 ���>yŪ�1J��I�_ס֧\���e���LYcP 4��N���l���-47�'౒}��g);A�E��'��PfX�Y$T|�0 �0,^��8K���r5�L�(��r뺸`ݖ�U��k�2�@*2q�j�	�}q�M�DX���Rw�U61��D�"�=	��T*�,��	��ϪXlr����zo?w��7w͕
��с]�t��PDO�/�ָ���҅ϖ��<�K�|�� W}�h�E!f�sr�c�NA�w�4[�v���k�`�f]]};|Mrf�ۅ�2q"=b����_����L��C���֊`��&'�]J����H�20���D��*1e5u��/ĶZ1pf���6�jd���-�_IU��<�C1�3��Y��0���A���!��u_�6���ߔ#�"1�x�FH�*N��R�'��9��`[��^����r0<��M�'�N�=���??q�pX��Vl���Uu���Cw2Y4Ƽ����䎮h�ԉ�F�)����cR�0���:���;(0x��<?��/��Y�lvb�:�$�x�V�:1C�1�sgX!hR�q�7��?R����Jd\y;ai���쌴���?G��(�ׂ]�ai�}���(���P	�f�g� �N�p܌0���+���͸2	��a]��d�����m�s�F,����|�*e�n�Z 3VMot�����A�;G
i'�[(��fߚ�{�h�!A�����w՟�3S��!y��)�9E�l�L��p�Ūi����l���ع͵ˉ
�q?b���/�_<��'dXݐ�^J�$?L�L,������!
^;iʥ3��m�t�5���3���V�\�c�V��9a�<lL�RFצG��u�+���k������Y���*�j_<D2��`�򊿺��t��F��J�uj&��bM��9oj1�E��]*9�.OY0~}Vm=��U��ʾF����~�6��^SY���<�\A��]�jp��C�^`���&�  x�j������0TУ�0�Q�Ƃ�<��|mߘ���6�|;��eƖ.G����P+Y�9\av� �g�8�ΐ���B��׮DqZ�c��fYqX�B�������x:��όRV"G,�И�|eR�ziK�!M�Z1rn��&��TBR������mg齘� Y1@�����e�4Ṏ0���V�urj��zg�"<ʓ1,���Z2�u´��o���aJ�Լ�L@��	=Ѥ���ƃ�5B�tM��G�z�5�8����c�2
�j6�!5�u���e��g�:rRΉ�9�V��u���A�����R���՝�t
����|2�"��f���|ЎH�.l-.�}n�S�}�������'�y�������'! ��-��_x)�����3:R�=��{f�֣�W�{�����<R��O�&o��Ū�a_��POe:�� �w������{u�{�9c$��1D�eq=e�uW�-1�ٳ0�~k�V���%�(��E�<�2�����I~�>�M�j �AiX)��w�7Z���zו�����q5�$FƩ�'9�tٽA�`ɗwDRW�+���No��B!a� n�>i+z��gu�nL��I�/n���*��y����R¬��uq����}����e�f��>���m��wx�tO�R@���U�t�iD��=����J
�ԫߛZkو��j����5�i���ƨD�d�R�~�^Z#��V؁-�������XGǩY�"��a�u���W
 ��L8�2t�@�M��zd绩�<<�Tf��HW��ߩ�^���-�I���zK�M�ug̎_���a���Z�E(��%���Ј\i?چc����6�ñ��^�c!�:jr�Ev���"e_��O6t[C��TSm��Or���ۊ[\yƗS��=*]�����B����g���"���re�h>�m<�[.N�<k�������Қ�N�����z7Pz��I�_����H�*�5���������@���7�s�KJBUx^?-�k��Ϙ4AҎD`�$
��܀�c�G|߰��3�Y�� �X��'��ܡ�ZI�y�����@Z%�AwV�����w!�!��NM�؛\�O�����\��;�����=�	��"�h�'-��ļW��[ ��H�&|��l�S�1*-��*�!>*���+2+���}2u�Z��f��;�
|@8O�p�<Z��hO��5�Y��h�4<�i��o�;��&��������<,6,�#�*B�����S�hʁ\t�j���f��T��QG0�b��2�'F�f������Z1̥>$�(g�,1x���w���_]�����q!?��1t@�ޠP�rs7�_�����k�w���*ϭ{�9��k4��Dà��O��*�����v�1�LW:#m|qME�dϥJ0/&,�<�r����?6��������C#�@u'dWm�)/=z�@:j�]����%���UڸAEc������7�)���V�0¦�1n#�P�x���Ep������c���CJA���Is1�~�����R�\(C��K�������%	kE�G8�[�zg7�2]bN��l�����wC( ���|���&�����a��Q����?fE�+�1��cpD����=u������1��`�����8p�83�l(4��̡�a��]�����c^B�<���$����,��{�+��E� �z�ԟѱ(��^��8��ݗ�P�0Eǁ��k�jaB��Nr��W�a�]�	�-��Q���6	g����'���"醊^���j������R�u��e~���E��3w��ϛ�5=�Rݙ!���T�LI<���^}���,z33�⋮��0&��M����lF�p��G9�>�̫��B�x>��HB�^DN�����&kr9v��C�]�I����öR$B��yʑiGs<�Զ�P���H!娒��8����|F����E7��;�)9+���"�<;��B$ �l��jdR������$���)���I��=��* ހ�5��?.��,���&<\2��Fm�}>˹�xS�F�I9?�ZՄ��PZȍ�)9�w�X[� ;71��(N!Ҧ��R����� m����~���\^��m��zt�'��ip��8�o0n�mQ�������6,��Ԉ���2ՒfZ�t �Z����e1,(L*i���ӻ1�9R*�c5�Q=�^b�;p�G^�1��'�:􆌔�\��4B0��[g"��^;)�Y�Z��Ġ%5�z��B�ǌ���-԰*Sp��`u|P@���AY&tg�I+�t�s�(3پ�N��]�a�7}�͹j���&>�堙=[�ë&#M_�V���;��^��(w��u�N���u��T��J~��tJ����7I��2�RL����\��!ҬQw�Y���r^�v�F���@��v��`�~���P���O/�m����
H���)�1��.����]��T�^�?��a��52�"�E�'@�C�i��eWp�S%G�"P��HoY��3����7���:}�yb��v���9}��u�ݚ���x��&��0�0�@@ߘ[��c%��7�j'���!�g�l����+���U�(����&}�zĈ����~�sU?�I��c�Q��|9�\=b�U�}Y>����.E(��*"�z�?ɼ�$҉]� ���>��*[�m�{���a���Z���BB;q��>�����=u������"e�.������F�׷��@�?��IF>B�T[Z��bs�A�#ժ��\��(�d~f%9mYe��Ӗ���>�d�dIH�C�iee��wnZG76r$jm�@���b��@�j��䅟�Y�&i@a��'l��A<�t23�&
4] _�z���B��)���L+~�	��WM�2'Uu��G���ŘwP|�PP��<��Y#�A��#4V�C���Y�����	}0nF�z��.Z0���R_��<��,��`���h�"&�<�Ce.��h�G�T�N��a~h�C�� x?T��O�|ṡX���N�o]��D����n �d��u�p��Zʭ�p+�w'�M�sΧ^�G��o�*j�`���|�'Kk�>�a�#�`V�|�i�2=�z����6٧�8���"Ri�M�G��}���gOS���OdV\�˾��;�+�gp��i?Q@Lap�3Y����Q�S��JN�=�c���fT}�%,��>d���[��	�Ɇ؝�ӻtxY���;���X��3��O7����7?�c��J)��$B�b��O2�9�i�)D}����Ͻ�m�1C�?�7�=	W�9#���'kґ�˕��:A��'��)�?�v|��!ʳ�$ɦ�J�`��bA (w��w@��\��o�(k~��mn�.+{�UZ�tI�n��pv�����5�83��9`���+�Ix?��y߀���PT�cI]��q����F����pũcz$	�u��V�!W�6l��y~-� {(	����n�M��XOL� ��r��1T��-�H�|����q|e���jh�KS�������$l4�5��:E���U����2w:�� �?̒�VaBG�;�]��j��Ccr�p�!��ĉ��Q�v�����Px�����c	�Q62����[ر�+��\}���me^�0�(��^��C�Y��I���e�D"+&�Jn]^�!�LF�ݩ�����GQ�C4�oM��*7P�P�8Lx�i�����Ҹ�2���%�	�8�U�K�q<:��8�n֨ޚRP�_��˻�ߪ(ë�����o�;tEC��_������}�s��!�>ݼ�#b��v��,�.c�^�	�Q'�aW7���$k�VCM�&�[W{�����4��Fm�zҦ�|w#�O9�?$�w�w=!Y��ts�EұΜ5Je��M�O���Yd�+�_J��f6�]N+=��3����Z�+]��>� B6���q�1�_�Qg k�F��;��:�����Ôj��6m�\$֍�2��gk���[E������j����b�����tC�Ŵ��R*�+�T��Ur"í�ɖ�d�Ό�T����kH�f7lָ�N�V
��ɩ��>픳6�,z�V@�r�avl!���q?'��
�qW��!�k�2ƒSq��c�Jv(C(��&#���I�x�C�M�9s�"R{u�ny�@����qي ��Qu*��鋼2�M���*à�V����4��ͲK3Y���o��������x���0j#���@G!8�U?�dX�_yZq�1#�=�b�K7ޓ�R�%�s:ݺюb ��Y���M%�_��c�6ycn˱��}�<�}C����33�,À�ι��!���mbP��xD��ɜ���!��>b�ܹ�3>�Ƕ�;�t��@6bh��}���%|����t7E��Ȅ4�y�6T�K�5\�����K^�� �U�nN�fc2vM���Z�	_��e�#�}�G5r�H���I��.,�F��j�>�Ԏ���dP$�5�&���K��o���6���[�-����jLX��E�΂�Q���6&*���:��D�^�cAܦ�72}��,�������d���u Z�uɧ}�NP|�*��l7~��e��J��HHW��)iw�����	��n�~�I�6o��:��׎�%����pqr��}t+RX��,p�����=FkN�eE��\k�{�b�:̩� �i3FN�T lG��^M\ɥ��>Wz[{��;[}�W���U�=�kG��Ih�M��u��t�����[cF��$�sz��N�9j4hny��ԵMل���`,��i��~�?Am�XV��|��jY§����i�N ������r.B�3�W��" �u(B��
��4��u����H6��q��e�{p�4
X�������i�!Q��|v�R�G�-�\�v��P��	R1M�K�ae�[�C��+��i{𗗫���v��`�?Xc�I�������6�󫂃SR�d��ua~I*���O}�男y�K�dI��E~I/�\e�ƃQ��/Ώc�J3��N*p=�� B�/P�[��ٳ{��IWz@��{y8ݖ��x#x疹[c|oB{�~r?��H_) ����"�n{e���KsS����@��y�����x*����g�)��M���(g��%鞱^M,�k�����a����~;�\�(n1��S�Je/��A���z]F+@�ƶ�����'�<S��[]p�tG��F�����o.Znr�Y~�$��w|�6��B��k��Я����|�hI�x➐��`1�0�^Rx�ēG������nr�i�W� L�;��[�g��6�����f���}ޘY�������Ϯ	 Ftn.1-0�8.,�x�Vv�UqU�ۃw~1:�e�e>=�9�q�۔֘JÓI�{���-9����o
$�ڈ��(������[P��F<@���9�N��Ɋ$k⊺�9T*��+�f`�&�\ŏ=2Cf��,�[B��c=�YD�C�N\d��ŝ�]u\�E5�,�-.Ǡ�]�(��[[k�ED���>ߘ��3&�����9"#xd-���Z��ɄF�JM'������_|����w����\�~G���\�B�b=��$�=�K���}��r&ȆZ���$���p����W�=�������/b�W{�j\�k%$����R�4�W�#�<k�	)����jEoFp��P�'�p�oiL�YgYE~��٬��փ4��|���n��}�d,��TQ7�00}����?������3����t3=N�O�f�[8aiV�]�+u�aB��n�rZ.`�v����r����h˳f�="�ZC�8�rp=��͎�H�C�p]G�f$��� ]
�`t��I�Ɋ��iVEh�.3���#�r��H�]�t	)�y���{�*엹r	�`�[fm[�{z�ǌi�88��覡%���.���+᙮��)T�>%�^h���)���bj<N�1�:��&�>{�߉�?�6��c��CD,��R�;䝒����ei�*�+��^X�#�;��j�'fp�~���B�d���2r*������J*�u�z+��@��5�5Fr�V%��"��}�\��
�Y�~�#]���T���FRPd}�u�V��ʂ,����ܙH�箂v9@��;�Z�c��{a�|s���b���J
��\�jRc
��_\B�l����3��-���\�|����a�s,:!@�3���<�ˊ��
H�t��L�$EU��� Ş�_Y��z����k��R2�t~)1�9�_|M�s>��)�]\�,�	��!����C{Yj�?�i�4ϓ"^]�^�iRpXK",[�3>MN��
�	3�a�B���\"9�p�B,_U� Y�c��
�m#�㕵�L�؈cX�?v��~\�Zq�Y��$RJ?1��\�<�i%A��t?��!�X޵�H}@������-�ﷁ����	���掲���I>k�3�@z/j-�WƘO�k�_��l=�U;�Jv�?���L�qտZ��� �Esp������l��9���4���X!�����AM���6�bj9*�N�����DmO��� ���@ٿ�b����QJ��]P�	���M�/�7#���D�MO�83�)�dlOG�V!�γ ������h��7G8{�f�[�v[Ѕ���eq/�3���B"*��!��Z���fMz�q,L	&�t{I�~���v�X�����f��I�¼&�F���Ɛ�WM���H�H�K�����@P̖(����9���R��J��oM얯�o����U0��[{������a(�h���#~./ȴ]�&�� �]a~|$�]�J$ߞ! -L;n*P\��1����uI:0Kb}����'��y͇.��V�5˕{�Uo�1�
�CgAa&3_r�U�݌x� ���9Yy8#�`*��y}'���<tGӼBe�;,dd�"W䌟����R��jщu�d8̒�pB��=�b[��1�s��m$���֟���b[���&)r*�D���P9B�ñ���3/�Bf>�~�ţ�����|8u�-���dް���E��SȂ���Vb7O����'/����)n)�RgNR9�8��q�'����������!h���&��ޙ�)V��QG�C�`u�&Ab����]sK��jO��m�Y��]��$��K�14�G����j�H��o��1��R���c4Y��,���k���'8����������L��?��Sm�5�`WRU�;U$��,+��"a ��ҎwL֫�?٦�:ZέI-�*���C@d��:��G��#���e�)ML=-y�s�X[~7�����YAo=����BW��A���¨�C�b<~�y���:q2�Y�Cy0Q2����>F�����"LP���g�
4Gܻp�1��yL%���}���C�y5�gz�ך��{�����
L����^)&a��I�e����I� |򆤜
�y���z�Q�(!��v�����ĝ����d�t�q���I����w��R�r����������i-�^�{���]�=.*c�[A-�������gvH|��~���fR�ο�,��6��(��P��\3#<�_[���P�\	M�P�2��S���$\��#$�+0�ͻ�玕_#7��s�,�x�][	\�>#��mߎn�526�EW �'�(�T����:U�1��&������Kq�[���]k����9`�Ʈ�y������M���,&��o��"{���N�}������[A�I���ؿ7��!����/�;`;�]~<ĥ�z�=��.X˵�A����{m������Ӱ@�����8)W �P��DG�N�hK�m#��w�+�d���M�Nt؞q�<L�I�&Q�95+o���:|W6?�kc����
���Vo�mg����";��$� W��ð���]N=4�;�r�Z�c9�����X���b����%ߙp�aP�b
�g�ϼu+[�C�e�Y3�JA�)SuF��\=����t���io�BA�:Sŧ��-�
X�KyC�g�s����sf�ʹ�+���܁�srz^x�>F�^m�X�bE���=�ٗ���X�yk�6GUⅫ�i�����k�xcD�|��F��%y@�3��eI������s�xD�Ԇ� ��P�Q�;�$��������W�~1��kxӷ_$i�SКZ�4m7���(9�o/H!��%싣ؔ�]��k���M���:䘖��H�� �
��5Y��N���.��P��砾�L1w����3���{����jQ��kh/ez�#���)9#4,��!'�n�1�����7��+��M�v�=������,��㚬dn�|�!D����=^�uФa�Q�W?r��<��#�:ݙ�d/�|����S`0+�2���}�%��R�}�J��?��˺�����";��fQ��y%@�_�0@0d�P��"2��I��0���VD�cH�j��h�.9��<�Gb��6"g�
=eD��0T���F�8D�.ϯ6�;z����*_��#��:)?�9W���K�m����c�*Q=�[i�Nٜh.!�J:o��ę���j��C�z�j�{.���������Go4	mћ�[��e�a����b�#���U��;E�7��M���hi���i����8]3�F	yѺ��YC5d��ڎ��0�g2k�����ڶ��6���`���g����#.ى��pa��M�j���;
,7E�0���Ѝ��Qg�x���d�r�/��5���X"M�sKg�b���_�:q=�5T��;&}j�������v*�U�U�t�"-f�@n�d.�wߢ-�ߑ�Z������C$Yݛ�2�3fc92nw1<@�m^g�h�vgLO;��vO\2�"�}����E�M�QV�_޺���C����誻��N��|����4��o�{��Z<!�`�#O�R��(�,�����Q�ST�,���v�Br޺HM�3iv�L��HR�!I<��@�q���G4�{W���G�Djk���+_E���:��g��� ���1g;@�s{�9�I�tg�v�l5��P��Yn¢�(�?y
��s�z��M�Cl����Kz#riX��Zf�#�o�d��X���#_-���Csղ��g R�̅�S$L��
*ӹ�;�^�2'V8ղ�m@��]�P7m��u��:���Uf�P�\���Rj��WIoN�uH�X���5�^��~p*�Ww!?��K�m�/�"v�Q>�6c��8�N���iu�Zx'��K�@[$Ī .�z�ZRayi(I~����tN��5!W��O`�NR�䚐���󓰼�����K���.^�V
���NO1�eB1[)
3��8T�Sn�lw}��� �1i0�E;޶�ىs�
r��M�jɬ%��,����*��l�x�k�?�0���hꎄ
�M�c~��_�cD��US����SY�|>�7n�e��V�kǹ�ؗ���Qb��d�����҇gS�d�A�1��0��Rk0K��^"�|�����0�<���}Z�f�Nd�ղ��~�H�
$S��K����`���"\�"lOޟ7 +pI4�H�X��r1*�|"z[��B�uq5���މְ0}����I��Z�
���H���y�Wo�J�E��,[�w�Y��u�1ߨqi��@H8j�<k�7Fp��TZx�w�q
�Q�E�\b�қ��t,x^v�y���ӛ���/���Jd�ɀ��HQ��ӥ$#
/��2��n���y�`��z�����x�(��G��7f�Ւ��x^�"�Xl_Y��%?+cɛ,n*,��)Ұ�2��S�GK��5�D�6E5h�]������Dz����?�B�A6���@/��p��5�D�i
|4��]��Fl��,���}b�+�L��ȥ��-"_8pp���Ԓ��k�\rL�%ڿ&l>����bƋ��aGQ�_f�J�{����w'�=6u�*������%�,��:gdm��{:�v[�o-woƙ5A���&���;�_���g�X,`x+e`������}}�*�դ��#'<K��x�^�K
Bi5�f�@���ὖ�����!����� ��iBo�W&*�u��#/j�ѻGE71���sSn�@�����@*K����*��7�CWG{�d�T�!��yb��ff���q�ߘv�f��!�wRm�Xw��y�R���"�Yy�,L��A
�1[���,�^�W� |��c��JA�d��Y_φ���K�����z�����A��t[%�?X787����PU?}" V{c��t^Z%�a�ז��As)�po����,h��rצ�NJu@����M��P��ܿ5gj�n�#�\(�K���0e:{g�ͭ������y6Wϯ���D�1#����3C�i�؟�nhF]���Uրz\?�|*�P��!�f�#�ե��vi_Ȑ�b�f��,���}~��Q\�g�\Gt�\$��H*����.K�`v$��n�]c�]�5������E���XK����_da�ޗ��[�$�*��s�&-��T	lD�Q�4q��7���^2��c�d�1�>y]�5�ŭhtzN᧘���/�/��Oa�,�9j
$�Sz�ǂ�~����u��V],��������z	��_�6�IMvSz�ޭ�]ˋ���
pprf��Y�b1#vK=L=�:�{��%�'��ǵ���Tmzچ��-ʄF����X���"�Yh	ŀ�L^П�O8�����VY��3�Еe=]ue/�tdZ�Μrc�^(Л�dvr� w.�o�hH>:�M�Bc��!Edߔ�v��nPxl���[`�A����\ u,8>H�ƦdJ+El' �3�md����=Y�vZ����?��T�o����m���Z��p/��c���x>z�~56��uwᴧ�*��+=̶� �75�.��bZb	�l,&���� =9Ϣ"X�Ux{7�>���y�;�| ��Y��˒�̮j0+B�����47)�oĄ�y�D.�7 ;�:G��k�kz�[�O���9�޹��b� ���%
,a]��to��J]�#��O>%W*���p:1<�|�<�!F�����s�T�:�|N�ڲ��{"�7&�*���{�
�-�U`Q+'y�a%6-� ��� �6#����k\�;�H�|�t@��"�($�9ߵa����QlW��,��9fPZ��`�=\pC�{"��ƐuSuԫhe7�K��Ԩ��������K!��e7��L<.b�2'��9oY��"�\��ъM�L��JfGQ$FBb��х����������2�<%�%)�w��8̾
�������s0¼S~�#�%@��9N)��[Y#7�i��N_s��l��F�󙪏t�B����`9���ܝ��R�D�*�����f@P�%���U1!KlX[4;�������w���~a�b��H��@(x0n�۳��@px���T�Rȹ��亇 �ϑ�����.�<��j�!��Xη㸬�k=~@qx�F�A��녩�J6ʆ��/u���	�Ef�����h� Rڜ��[R��ڹ�"hl.���',�[�iNTi��	xY|nڸB�j4���Y�V��3���p�����M��ߑQS��3:~�
:�Q�PY�Xnx[�� ��n�������1�`�N��x?���e-^cg�<.�Z��C)�I�-F��.�S�څў���~ǆ�6�5���c�����!���̊HQ]��c�M��W�%*���|�@˂�j&/"t^�=�����Z��hbo�cWQ|C��%h���5�)�XK�	��G���s/�Yō?y��sx��P�KjGX�t�S�c��c��Y2��(��LF����mpQ��~j.��E��3�:��/]��a'��4:h9O���Ӫ�&[D�da�#)�r0���-M����.�>��A��u3�*F���r�>�,��m
��4/V�H�O���������GZ�U�cL�\���ۧ}g������,�5��x��Rr!H`��]`��8�ON�"fvݻ������Ϲ�5�kQ�NE�`�Dn[-�0��F����U曀A��KHpW _����[��`SO�a:�I���Q���$�u�E��*�i��O�-jU�Nt;`�;��|(}y^>G���>���@�~\/�_�Ob��k"��h $Z��e�9��vI3�ã���0X��P,>B�S���<R�a��. �����Æq$^�j+Kd�aH�%u��(�z���1��b���ʁ�u	��� �����;N|M��ˡN!^0��O˿=P�01�G�4�+a)<����D��!��#���6=e�אof��l�8�䞑��|���^��-��l,1s!.uE����\2іE���_�R#F� ����fwG��\��ol�ܐ*X��ۢ�.�c��?��5��q��s�m��5񑳠X+��wɜM-�dM����g�6�>��Nl��g����)�Zl��_w6�qO��ŶH�f�vx(X����6�ڽ�uJS��XE�\L[¿R5�:zc��/f��3�?��w#�y�O�!���J|�&�
�:p�����"F���<�;�_f$pBysR�n�3�P�)q����d���K`[W8[� ()��7�م/M�*iZC_�0��Q��",�UD�P��&��p�Н6��7�p1�j���=T�O��y��ZN�:��_�8H�l[F<�����K+_:&��v^|��3O��;KTz$�Z�n ��O�%������v��s�&�`�e�e�z��[Vy����}�����QEf\��]���9y�7���{lj��A4�L&1�j�n�}m��al��w<�50Me�@�u�B�ɵA��-�n���b`�!r��p�Ԡ�)a���#���3�xƬ�kș��CBϛl-��>,��Mڨg&�-���$��bN�l�9[��G%���L�94ln@s�o��ӯ������L0�,���rbU"?�Nz������H�']IQd{��ɮ�2s��67�#�3�{ݹ�a���'�jE�kN�{��_<�����v��XU������� l3$��qq~�xc^4�w3����9��^Io(b�]�%�C�����U�opQ.�IL���S�,QX�q�ȮB�GACR�Er�ܴ��)�g���y�d�����T�6�;Z��3S}HQi'H�C*G�%7�8�Sǣ�2�_zx��r�)6��Cl�k�h$.�Q���jP�V��s��kF�ؿ*h4 j��'��D�F��͔��0Wk@:��K��;�ab)�2I[4�#�%q��r�5���H���&aF�y���K4i�0�]�t��O���zm��6��h]c�M�q*/[	dʉN�������2�貝�| �o�QG��>绍Y3��j���hg ��G�rHu���c����#�����~q�>d9?�V��M5dw���b���Ħo��SA�^��c~���{ j��S�h�</�#�F�0�a��i^~���5eO�A]E�o����m(�9f�j򊐦��%��g�l�-��<8X%�l@m(�QӫڟV����鮏+2�(7+I�K��"K[��+�{V��P���G}��Ss�Uz��[.?Ǻm5r�f�`�X@�h�ө2�e�6;{'�E�.��`-l����Cm2�����y����щ�ۅ-��#ט�\�����t�B�ԣM�tm�wۋ�l�8s������D�G:U�,�������	�KLsZ�Ҍ(�y�� �����]��j����VB1��B$D\Ge!a�)��r�yF�,/�as`�X�(W�����M��i��ѳ���i`�n���]�%���Ǎ���aQ����X�k8a-,j"VȘ�Sf������X|�@;�M	z�5�p�Ck>���0$����vF���o�
�L� ҕ<6��� ���]���\�d�3w/J(�� \,����jC��\����`�[�FLk`�z$�8��ſŞ] WU��8��EZ�"��fج�sT\�O�����)�Yb�Nw���sB8E��Qt���?�Փ�f����U��:"�ճ��<��%N����Ҧ&}���7�O�CO��|M���Fhg�YQ[x�A�	�;d|,TI婗�CO��+V@U���=:G⾪���#`���[E]7�r�w����tR/
Q��l1�6��������I�{���۩&�꼇������')��d��wS��T�Цs��ee�Ц��
�M�S*Q�/^USk:�tc��P����e�$���RjV�bk�SQ5v b�b<����X�	�A]�F��Z4�ZQ̓{��n�@�̧�$���v�	�����(̤V,�D�6v06��$wqsl���Y	N���+���+{7����߸c�0y>�G��Y�*�
�!�Tu�\<g�{���MEKI�ч��ʰ�T�,�_���f�~�ʐ�'FV��}��=����4��vqoe��+��\��TVg68Y��?��^nr�� �����?Я��CS)��Ԙq�<Z�D�~�����y�QE�~�6>��֠�推uBGEE�0�`F��L�)TO<u0[��$�����	A�4�.��)��IT2�'a>�����,y��4�.7�_�a�FCl�_����� -H�p�b�/�O����D�?�����Q���?��ᡱ�o_�z�m�c楊/��v�>�:�ݿ���a�[�7���਒�Ԑ	x�@��k\H�T(ާ&+$(vdπ�3]{j�����*.MN�4*�f<�wS`a���&;�
