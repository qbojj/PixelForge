��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����P�^�Mqap)%t�?�&�Z�K�*���~O��in�ÇZ2���RG����R����k:�H���QNOR| ^{Ua��M��m�:�$���/�s�~J{]���Nh7�_8���H^����bu��<H%�m�i�9c&*>�5�Gd�6ΎD�I�#�%A��#�Xq!��n�����"WGE��P�0�£�T�	����H.�6�P�W��G���DN$�q�`�S2��SňJ☔+��ʗ���{f�$��Qp����i��s�h?�������-5y�Z�W>��/N#��)#..���7�t���;�\v���fys�����n���s}뛨�*d��PEz�V��I[�x1m�*�"�����47#7y���eU�g��W��*��:}�ۄy\���ߌ��ɺB�zg[�Rՙ�e�n��ʢ��Ŝ�._A�{��+l����O��~=`�e(�&���3���]�|�QlD������u��DK*C��M�;���3KNm�����~�1�&���Ҝ@�W��֦!���n0(7}:�=c��N��ŷ`�9�c1�ϡ�^�+��_&�7Y��[ؤ;,tX��_�����U��qn�Η/�P�4�- ��^@v�b�����ZU�j�#�t[�Ҝ�j�̐/�Z�Į��t�RL��)�W�S-�|&qbu�Xd��l���ʧ�~W�j�R#��ɑX.���LϗЪ�cBX"��4_3X>:'���`u�Z}�U�fHdLqd�O�������ЩL,��o��f��Y�XQq��W�60��j6�@ВI�
1��A���3��S%dj��a�3��8:������rS�p�����_V�W��GR�7r����֤͜J^1F��}�/�b-���=��gP��O���^u��SV=�`��$�A tt�=y�I�im���������d&�&��2�.Ɗ�:�o.�U�nw�߱�/9��b�3����]���$t�s�[B�u��
;������fMw)�@��'�)m��-ԶQK>
�}Z�H�'��'"��LZ/;���b1�AĐ)�
E|�>����U�������{?��P�,_�q��e�$�Jg�����W����6���+�a��E�0�0�+��~�8\k��t�n�p����̓6�d���{�k���n��S�3�>�U1�����Ib��eG��{�Q�����C���~��[\�l2���zt���}N�ǘ�J^qڙ��M�|Y��͖)(��9f�0��i>}���kE����y��ص�k�./k��no��^��U��k��tF��rhPE�?�H�k/S�m3Aέ�?1��^��z��6
���
���#��GZ�ʟM�̓Z�I����n��Y�!��������֎6�k�j�ӗ(Q�Y{���#�[[�ڮ��⤙��^1p��A�yW����v�h'zӺ���P8m'�k��W@�z���ȐYVxQ��V4o��zT��\ Df��]���аtS�P��2E��~@�+�B#k��B���P�kr�����@�i z�6QX���|2�k �!�`���p9�l�VX����H�ҾMI��;�w�~���!�������	1�����p�.��@ʳЪ������cZ�1����48�Ix� ����>q4�\����Ƴ���T(�a�b dH2���>�J��vǰq�|'e��ҧm�/��q�����	�R�y�>V��6y��?�R�j�3���C�^S�bj�^��1�4���v����J^m���xk�����B�n:k,��n\�V����K����l~�Q�u�G����~AI�fa�X�3EET����7_���ͯ���|ŲH����+L���l�~�Ԩc3�CH�u��0���}�MaT� F�*q�ϛ��s�ސ����晞�j���5��d$ט$��8 (O���֜�:x#Y�Q�P��f�[pxH��Q���(B�7Y���#T(�L�5��|��.���r�f��ߖ7�B
8�P��cY�nBR��I�/:=n�Ν^}��'�6���H�N7]�yT�:v��^ӎXIl��^�SIʘmK����d�yVuK�+���v#*f뛾}۷�r
$,.p�0�ۘ��a����h��UK9��ْ�l�r�s���C8¤��? �.��<�iQZ�TH�I�y|I��]"���ghD	����*�=|.�o���a����]�����B�b�R��hM�rlјهe@��U��h���׃�-�"Գ��~b��T��2h��mo�Jz�DA㽠u�5��Ҩ�>��p��ܾ3;��+��O�ґ0�۽ k"E���
Q�P]��D|�񚻱j��D�٣�1�f_��p�*��7�\L�_7��N5F���m�nm/��4�����h
���7q�\�H��nDQV��و�<�^s�@UVQ�B��[(�˹��p�ܹ*�e��ٳ
<ǔY��dU,�aƦ��s}�P#*T��p�/�����wC!�3�r����1�~(g�j뭚�W��U}L; ���9�k������Ԃ3��^5��"h���.Q�Q�xqq�%b�"@�]9����v�R$�*l�3t� J�%`M��Zo(W1��^ly�yjg\l#�N��+/�2�ޭ�j�;�W�&[�����+�c �m1P����2k���dZ�	ƣ�ρAP��p+�,M��Fq� e��� J�q�����N�S�l���Pd\�چ�D��}X���;P���~cg �Iӽġ�h�T�U�=(�rф�������KW�Ԅ�=���3��,Z^��P��c�1�1�4:m(Y�>��ȪR�3�P���{��*n�6��㟟��ˣ�QNt9�V`?box�bc�aݻ��K�������@_O�w���Ԑ[�$�.N>-��V<��T�����⌋뒮�#��8�Mή;e%����>�2���XǠ�.�{g�@��Sfq���s�h�?��!]�~���zn8^�S��,�T)�bE�-��b����	�%a�v0zew~u��.�䗦�&��m؇n�TN�������O���
(����M��������JT��;R,�\�Jʠ�9J�(~ʎ�R�:'�Z�KdJ���
	�r(�I�@��Ȧ7?�l�s�n~p�s ,�/V�&�m3Ȋm�lt��̐�_J�3�QyL�i2�g/�����H�����|����������Ѵ<�% �HW�l%�s��[�<Cp�%|�-�@�3:�҂�szb
�WTH��N��~-��S�f�ֆ��&�^���6���:�u^F�خ����|Š<4�}��Pn�H��g�&+��VX���������:�@AT�G9Zo�Q���4Ž��9�Y����#pT�d= ��QJ2*y��B�T�ZD�Qzx�Zxx����!4��5_?����������C��D�Dɋ+h�a#i���^����,9������jS��Qr��̑�<&��H�o/=X��+&�C!��������#��J�W������V����L��I��vem����gU��A/�6N����޳"���<���IT�]=���`N�CX����_�}*s�W�D��V�U��r���DMk��hP^Jk�I��Ҹ%B8�f���C�l!���U���сk20�/��u�X��9K����2��;3}�Y��%G���	�'F������G��{�浮��>��B��j��O��4�׵c�-���������T(S��ZY��[�C��t�סZ:�v.�;��R2-D��V���>Z�|8�{i�,Ƭ+�Ȅ�C�&B?..�f�/�������q��j���M�嗱l�v{3t_m�� @�V���%Ӄ#8�#w�K�aND��7��iU܋߀L�j_򀩰�ʵ�Yd�S��$����K̛jbl����z�R�U.}�2Ԑ�-�z�y �s�K^�������1��KU��QI�����L���V�>��"���
E�.w�����ͤ��xvi!,J�l#1_DD�ʳ��R}�_=Aq ���������$՝y���4 �����рN3n�c���������~[OLa,fD�)��j� +��_y�xc7��zNǐ�_FY����T-f�L'g�/�>KH9�UA�z`9k�y��x�~ �����y�DXx�=)�&��Yڣ�C42�,r�.�r�3��E���'	�k~XH�&���=�G]BD���-���D���*���\w��zޛ�Z����7[݄_
��|9��2ӝ��$P���M�L�)�֟.ry�K@��8�@L��f1��Tc����Z(?F[l��Y3�������
N <���S��)s��?+M���|ͨ -.Ox�u	O�"���g�����c���&������1��7���,9�^�|�M�t���"�)�ɔG�.�%&�#ҫ~[��x���U�
�T�#��נ4�_������vt��0�7�-�/ �3'�r#���	P���E��OYVq�<��
8�����"?3���0u;ĔM��E���LxL.Ul�O�`��/t:H.�aVI`��iA���;��PT�>��(0p`�4���r��(:�����N ����t�P���Ɠ���~
Bo�p��(R
4�	[̞Ա�>ج����ܬNI�Z1�����r:��&�"������G#���
���	B�kJ7�L����-��G d~A���K?�)���`�H���b�ȥeR��FZ�<���T�S�]�eQj��߳�kyu�I�����ŷ�'a�J�A�i��L���^lsH3���������a�&*L�q��V��Rj�T���Y!�¥�5�.�j{�����:ϛK����� �sg��%Aol�a�f�򅶢C:��?ĉ�吿g������<��`�G�&��q��8����3fO�t��m��r��b
̚5����&.\�xH�0�K�,a�Bcl���
 ������{ȼw���w��}7�˳	!��!2�w��_�����e��,%�q#~�H����ܳ����� U��\O�����:[��p-vMQ�'6�,�D'�7]��=��yo�8j\?���#W_�{Ǝ ��g���e�~�LySu:�(�>'��z��r|t�>�w�IxoU�_ ��9�/F9m�x���o�$�	�$�N��?�o>v�;�05�麖�\⢆#BK�Y>$|m�A |�x�՝�����w�m�"ax�Lji<A"�(7M�1J�9i�Q��`m�'פ�t$l^L��!�� ���>.�S�U�&�RyЄ�(�7����.�لT`��2����yP����֢"$ΘV����6�S� ���t��LC��ĕ�O��M
F�Ϧ������Ja�"o{\���T�G���bm�l��}f � _V�)��u:�M�� �Rf]�E�1uf�-�7�����ɽ�[\��� v�:4O75�q@g�������1+����C*��̯��u�;�q�_9!�b���� ��vY ���\#��+m�{V�� L�M֪1tb���E�]ŃW��+gt���:F+�Ŕ���_t�̑4�JZ�Z����%�qrq�*i�ib��<��f�MkmZ����^�ٴ
�M;55G͕��xY7�L���㏶��!P�E��H�!G��&B`��~N�0��n��9�S�뾼=���݄�#�45 h?���d.�`
�?���E,�ۀI��_�.����Z,k"^�q����bݰS�etj6m9�۬��,�^��+�֜�~������r�V�;p@&\��������B�g:@�N�y �!�� ��khY,K��xB^�v�'��C`�k���`�hn��A�@{�n������QC3�\z�aC��C���J��)��?,!��$����tey�Y��xjb=,��xW U��D&��P+aP�S[�C0�h:���Q� Ȳҩ��Y<��f@����rQ�{=7��1��ܝ�󩇠z���j������G2���6
�fj
 ċ�X�u%'�����Ja\���XJ�cb�9�ga�6^������ �s�|��sV�z��=�)����D�XЙ�\Jt(�s~����K�E\r�ˌ^��H<n�\?W"�q]��xb���+F�,��]�%wQa�Vu�
v/ȁb_J��.�����L}=��/�L�>v's�8,�/�>��q<a���Jɐ�S��KQ���k:��ܶ �@�}�SEH��3�>GX7Ղe�~/\��9�I"���0�*���ٱ���U�O�m�9��Vm�2�V����F�ca�eR���:��rt�D�B1�y�K| �/�c��N2lIH*��_����h%��[A��t�c��;~��@�m�n5
�K	Le@�(;��z��&p���g�_߸嵗Y��*o����p`0m ��6��������TƗ}��G��r]MG�H�im�9��vMV�����#�y'�V�@x3">���4#Ū�ًGb�qwT��b���M�A�?if=�0���[�&��b�݇;�>M}'�b4Z�T��f34�]F�o��Cl(2�o�p���E���[o����p�Q�W�
5+"�<z�����^���Ry��߷B�?����t�y��j#kY�·S[��0K%�G7l#���SM����� ���}j%��~�����	}b�i|b-�YI	�W��P�F�m�����eC�C����̽��R�ghQi�e7)��-�?�2���͑y�s�*S����\&U!��P��˵�w�OQh��W����b�z�(띡���s;	���Vv�9S���6X_�2������/Ңy>p�\*Yv'���b~�{$QG_���
׋�dԷ�aӮ7ga�%:�4�ѧ��|�!̄�'=g���-,\����c�Y��RW�v�`D�`�]�{egɦ�:Fo?'v���t�75d����h��2Z�d��Hm���d���٫�`�����Wt�;�"v��90kůQ'��F�1m���~�_������f�2~����Wx&E��8{Fv��ҟJc*Qz�H��8�N4�-f�F��}f�j����3�z�FN�?Q��L=����p���� ��[d�f�� \ݳ0`1�^����W�=sI+/�ru�zdSi�#��t����4�93�E���|���3E��8WG�Ņ�-�hS�F���ፒ�,��V�9(��l��#K�����p=��/ ��%����|�9�z����h����D����j����}��H�D1� ��R?��ڞ>hV�����6�ǼVۜY����P������!\��ٷ�y���\�t#�M�s�s�� ̅��t�����"8dm��:��p"x�'i�z:|���&�&����&GqP�0R�*8t5J��l����&���бўU �p0V���4���w ��5���{����A���ۈ��٘Œ��ݐ���h�%$ʑ>~�2�H� �JU�����N�|��O�p�v��e���ݓ!+#�GNz~�J�@R6׼�}�8�}¸�N0�4������w��}yG!��$�y͊���T�25Bӕ��v'��|�-�4�)<ly��v'��j�c��w���P�{7�к����(jB��a��-�О�l����Gn�2�@'sS��3��}�	�+��D^tгDf�~V	�.mlA���#��>E�ӦWx�C�`��XS���"�i$��4�����~3��c�(v��]����� �o؊�'����f�Q�Nv�.��)���m������00c���;���7rR�Ǉ]ꐓ��gMh4,�����t�de'���"��.�����pa�vB�)I�}s:}>��-��f�N�e�w#��d؜)��@�v�p����\��h��p�%��.N��"����Wˉ��]@�E�\�TgMq 8�CR.}���=�<8z�zk"�>��C��JDp��jE�iNi4j0�*� ��e�n�^߻��	�^bq.�6�o�f���^o���Ɗ@�֡�{���|���y;����t��Cdg�� �3oϏ.r-��ח��&bR���~J��fSU���8m�0AL}�1]�����{7<����z�>�����@����8����Y&s������oE�����Xn�ۘ�^O�bBئyi4k�R�y;�~�zz�ǌ���$����W��A_~�:�`1��y��xԔ�#�r���ib�^�@}�B,���'kg|�*��z��j"_=sW�^5�WrX�E6��d8�3N��r8o�<o��'?�W�T�֐2��i�:���:���Q��K�O o*X�R�]Iv
�_���1j�R���&}����/���%��CXZ�Nњ��:�s��z���.���?�T�S��fz6��U�2�rpc�^�{���t�v����R�`�H{�[U�?�;sj�@�q�l$�cIʸ@wu�31º.�v��!�.-��lc�Ǌ�����5�ǑPEILPk|�����2�-��������nn�Q������E!�hX� �d��Hv�HG�ɻ�'�.��! &���y��ix3u�DTb�	���M^5Y����dZ���T�8� ʡ�)�����6puL���Ei�kي �7�������ri�@�(n���>++�ߊK{����?���7���6�k�J�*�l������;2�"�T�M�2m��h)�R����+�$��s��b<�Ҏ�y�J�x�OJ� ��GR�����dxT�r���~�ߓe{g��F&��aÕ3çQ:�.'�6����2�� 1�"�5#�Z�6��
,w���J�W�O���Z.E���1j�1��3R���)ERhI�RY�[��&�Z�T�So��B�T[erf�z�x�Q�W�EPm��j7�S�"Fͥ�j�{��V%���b;���=ܪ�n�Ű"���م�� ��7��H`3���.����}V4t��f ռ �����������%�臌�g��+Q�YFu������o��(\85x}�%
AX�2�1J�I�Q�71�:�eo)���Yt!���wE�]y@!����^�����Y��{])���H�Z���B���m�U�i1-��&4�j��H��>q�;*��KE@�1z���M~�4�k�YF�ٜ�W'�f5	l���h e=LT
��ym�[C"B��Dq8`+t_��,u�_�4������ ����r��#�e��E�׀|}@Q�"ߨ\�ı����Z,�� f�K�����C��=v�^k6VJ]�Mml�ā�Q/$��{���(r��/�ʿP���IC�a��ѭ�S��v�@�rq�>Atm�|c��\O7�Vnb��n�>Z#$�(v@%��y��=1=��%�~�cgW���ҷv��Ә�`�4J���p=�������I�xCÒ�R�����t<��o]�/��(��c������o޴�X�e3�ژ�5l�0�>��>U=�.����E3ۿr���%~,Lb8<��-p3^��-�n�V�}�w.�9��Vq��_��""j=����U�!���-��_,e�ڜ�Jq!cy�֛���$��2�n�M
Bm���Q���I
���)LlD�{L���؃�㰆v*�����$J�g�z�2��Y�g�K��ny/8ѲvavG�ʂč^�L�2b;qd�'�s~�S�]N� җz���z�|�H��f�qe�L,����+��b�T����>>w�e�z~C��d`��:�툣���6n���C�v��I+��?�c�t��D�K��N�{�T��n����+�����F�*��7B�;� g_5�Ӑ+а��m�xcv��`��8s���%��j�1P�W߃��j����H�ޝ$!�Y�#H��k��%��O�WU��B�zB��E)ш�h�	������ڑpy��ϔ�=�`����[+�����w�oM���T�Ԑ�&%z�4�͐P�t�2577n��wX~@ę ���3-:֗��Mf��ON+>J>�ޔz���Kd#�T�qZ3Y7c��9�� �� �`v�����zm�2?kW��X�|�"�T�N>���e�͜�$IP`.��]I7bly<��=�xl3.(�͉'���@�7�����!�\'-(�o5�xG�0���k޵{�ݏ"j��.X�ޓ��G�?����^��H��9���>�GK$2ը<Z���K!A�9�f�7�܍S���D��wX4�mQ���g/Qǘ�)NkvW4
w�H��Z�\�4]�W�)G%�LP
y�to~��xy�;����d�WQ��)C��i�s�*Ǆ/j�8vk/�v�s��0⿱��\�Gĕ�.S	��p
czd�Ћ{�bPF�{���阖zg����� ����lE����n�~�B��a=�E�qW:�1��Rc9Ž-�a�h���'�)��P��]h��Q�Tz��۝�k-+i�����-��$�P�_H����]\���^A
��b���
ib��[=Us\8̺fr�~���&Fׇ�(#���yTE*��5�3©Sf��+o���w�D���)ĢG�\��;_~by�2L�~���q/���=��UA`�c��[�pn�U���=�0\'F��&C�F���j6~�2�O[b�y�\��&��\�4��kdJ�BLK,p�a!��n����Ga��򴺪��{�T���(L�fez9�Qև@��B��i�����v�#/L�}�	�r'���1�%�#��Ɓ����V8���L)[7�V�!䗸���v���6�d���}���ة�V�F^%ά�������}9*�Y�m�w �����L���N[a�ϖ��q��l~'���_�E��3a�QڨJp�ԩ�+���4��"�����V�v߾V��h3�/�@ 	��bu�>��7�Yj[����6j_����38
=!��ՂR'_3to�X�o��ZH�G��Wȹ=-� ,<e�,�����H2�ˏ�cLAmm>=::��fʒvc�<�(D�N���N�F>.�Y���|�&pL�=4��aˀ�����aR�^a-�C$]���Њ���0\��C��p�,��aT����|^�7������~����7rb:h�0R%�S��$���,�WP��7A`��D\���S���Ut[pV�e�����P�:�!{�.g��Ѷ��<��ñ9�TH����PI�
�L�e���A�k�,�g�����`�s���{i�P��ҟ��D�&R��L�L��-�z��z�@������|� ����_�S,�G�N��q�U�S�d�л�Kc�j��3Ӣ���()n�CSi�k�8�h9�4r���^|FդһY�&G��z{�<[ޛ�{:E@��VH�%�*��?�*DϪ��7RC�۽Ty��"��wRJ���I9��Z%^.��}�t���6��m�.��*�Qo$�nK��c�4|ݬ��lk8��d���/�U2�����ʁ�K�bx���X9���~��BJ��D�E���$ ������ �5}0�ػ{qQN��3���l6&��bRpY��x��fW����nT�����1��cH=#+'"��7�7�[�\�
IV���;�ZT<~��i]$h]ӼB�Y��ڵ�sm�*f%šs�F���\����
i� ���Gee�Y�l.�"���T�:�j����P��ǢT�>� _4�� �,z���()��w���l���P�O�o<�2O�,Er~�1��zc������!��/Z�:J�a}��0R&�+������s�F��{��r"��:u�e�mE\Φ�<=]����%65�}-��q��tF��o�D�o0ľ��:�?҂'����ym�,�>���V�0����/��
�^3�~�����,���/wZ"?��1��PD���Z����$����c�F-�juMt�F6fk��F�(�
����ȥ�����#N�3�swx���s��SJ�~
����9p��xV�'�k�:�M�hw�Du���)'�����Z�����/�s�PL�{%�%���ԋ,�1�Y����<�㊔X��;`�p��}S�� ���xS�@�/a-������� �}4J��#w���`͉��z��\��2�v��E8:Z�O��T����[~yw\�6�G����Ɨ_�س���i'N�C6	W��/����s4|���'�b�68�)����%��Zl���N)@1|i��xb�t��й�
�}��uX	)�� �e� ���6�� ����C��pV�b5���XT��o�	�S��"�W!w���!⦄��O�Ar�H ��|	%3�:Ų��=k�7,�`��D/���LZ�)�Z �
k���L,��! K��[�8���xE,�B�H����ʝ���ɩ��Q���g��L�ԉY�.CJ��+H ���H& g*���G3�Bh�J�N �{@����_�˂�O������Ƌ ܪ�;ʱo�ܐ��Y�7�o��8J����5�'M��g.XXIh#���Y�A�d�IM��������6���Ғ��T��>b�Y�8��f� s�L�+L�����)�]RS�%��!Hq����os��g�N1�׋����om��;M��u�s:z�v�)���(�/y��%)����1 ԯNo�n欃�6�u�|Wz� �+;ѽ���SWz���I�ݦI��������?H���ia۟M�)}��L���l�W����tY��t�w���� ��5�FLH׵���<�l=\�p٠W��}dVw�����f!g��3����wZ���N���8�C��/�EaR�k�w�����(���a7��?3��x&�FΓbxK��ݑA��<�ue~1��iӍ-ҏ����B/=�*��:髍֦N���<�����P���G̓\�����Z�k'9�0���K���a�hc�Fl���=r��G7��j�x��2����e#�w��x�5U����"�P+����ܚ~>��6dS3T߁�M@6�u��qszPz�5�>��Hok_����\"�(^��ۿ�����{���z���Q�CxLd��=�4p����v��zT�3ݒ+ޜ�$���7`�n�/x;���3�԰T�DY:�����=�:�Ǟ�m�F����d�э	"�����xA��Ug0a(�G+�h�0q��ʈ�]���2k_A�K���Y�횧]�
������1�-fbL�i�3�"�\M�~aY��I�c)N�������|ĺ�ֱ�����ßLکcf:aT�=����s�봬��r�U��U�X4y����u��Y����Wb��*�������]��hദ ��m���/k�v&RF=#}�R:�B��Բ���H2�'�y{2_;���nL� �gP@�q2�D�����ߧʽ_��MF!C!��m����3���gUruky	��d,8Xp�8�*
��B��k�P��)A=�*GXn_���TI"�9�#�y���cx?���=����<��t��9j�� d��d����҃3n�Q�ݬ��'j��nM�9�/�w��22���3�I��>Rl4|0���ϒ-�9�ted��3�] ۶$�h`kV)��I���<+}?S�KX��;ml< �V����d��@�R�ʼ�Vը��*'��������)�_�^,Ӝ*h.��Y
�Eې�/����WI��
��	�t���8$~�yt�@��S��90	�������+�9�V�{���v~�F"|��\`��+��	���jz{�E�0�7m|B/�oٯ�Ix��XqQ�
�׬�h[@�yMi$!�wYEٞI�k�B���u	��9��=lB=�;o/��;64 �}��g�:�!�C�d �<�z��D
~?a���T�w�F�;L��66��_,�z��VhL��;��9(�`S1��%��d�*>�y��������̸���xGIٳr��|�hI
\�%�J�v.c���c���o���ᗋ�䮲U�+|?͟�?�t��6����%��]H�ff������9��	�+�h��m��*�6����o�i"[a�W�ad�ʶ�x:�A��}��x=^�+ǜ��xT��$��.;����;Z���dw�������y?�i��i1N֜fYEO+1 MS�A�&����]��〧ɬ�ؾL)~0>efʰI�b���ćq�%�:e*��zGf���3���r�yw����B78ռ9+��e�5V�����ª.E�L�D�H"p�t��b�|����&U �QфF[`��\�sJПS��A��63+@�6�D�>�y�%p�+E�UOU�2@1��$7���e]ű�4[t�k	h�L��V��>�wB	��t&���X۴a����4�`��Zt �����f���P��0�f~Rc`�����G%U�?-����3z~���s	�Ο�����s2$dD���)kf�&���-��q�Lb�,�hr6I���t}�+�z���Ɓ�6e@�a�^��J:�������pӆA�uL�+�r0�s^w;RR��3q�
2`��Fm�P�b�'x}'��!��L������:n浥w?ϋ�R�$:�[j(̠����<�n�S�_��<����s,h�G���P�[T���JgZ�K!�Lq-�c�P�wT�t���p�����]�u{��H�?���k�� uhMcpG=��b }�M3w�}ę|�ǲ]��z�G��DmI�C�}��uP`�,�w�E�^�wd��蔄�V-F\�Mdi��*<��e�\�޸�ڎ�u������b�(>��g�v��Hp���-ćM�E��>���
�%�봕<��r�M��4�4u�cy�%t�}��L�v+�r�3�*��=X_���%��C���y��w�
�)/�M�l`������O9�Ԩ����&Q=�=]����%N���;Tp������gI`�	#�؂k/{�0N�(�JPn�#Y�� ٮ���:����ϻ�^����X-B���11uj�� ���QZ��C)�Fo�!zhU���%W�
c�B�-'���9p��an�.fw pGbz�\ݿ�|�B4��������چk\��K���g��`wT5�W��Fi����	�k�y����E0oCy�.0�lsl��g0�NcԤ*c�=�k��^(ն�Q�+��6(ǍZ$��K�Z�,/'���>��Tht�1�q��JC?�;�J�=,��StP?��A�Z����bH��<>z]5*
}<��+�-9ڎ~r���e���L�D�ׯ�I�u�����k��O*�i�T�1���B���W�444z��yM�`���f�{���~�fC�c�@�o4趡��fs��΅s:�v��a�pt�SaS�k �$��/�8rf[q�.�K�d�f��kz �إ�/�\B��煨u����M�wu�r��o�G�5kF+��9�.e��WbX�5�'.%�q\7r�����RsB���� 
!D�AHm�ʲ����r|ң���SSR���#���ʘ��%��B���=]�9ra0�:e؆b�dݰ�S-������g�u�#�=3P^g�w�4h�\k���P���8�=�bk��Y�HJㄒs�%�B�5�����Pa�f+VU��+�	u�X(�8�skU��"�gĲk��:�u>�)��|��x@�e���������r)+A�M{l1b��>)�;������0�UDqTkL�33<t��/FR�%#��&�q�.(��Գ��(d3�}˕ݮ���a�3�s�3TP�Q��z�F?��jq�dR�>V�K��[a�>���L��dc95Z���f˘<V�cQ"��̟/90MIw��J��2a]4��+�:�E0r��V�U~">���]6����9�rGWF�g��^d>�{� �j�J+��f�]\�m)��c;uj��'Ǐ����Q)w�8	^��n"��A�� e�(V�'��v9�Kk���4pU~�'�.�Z��nM"��� �O�\_����7��"
X��8��Ȃ&zUl��)+�]�;�vg�9U��}A<쒼��Jv��멚�b&����PJ'o��Z�N�;wನH���s�7��$��v(Չx��a�\�)�[��Ur��`�0� wC4"����2|�)���������B�[��j��U�y�����%ս�5
^�-o!�;W�k�IRy�),v&6V�(�w��jgʩ(�w��	E��t�QY�E�+�h�Wב�2�EEO�,u���ܬo��}XO��?|�51��ʫ����ۯ���dJ�Q�jx��JH�_��K���ؔ��|X��Y*�I݁-K��ch��݁�㾳G1x0,�,`�����=��А���P�j�2r�ǭHzX�/�ta�1�?ѭl�]�H����d�	NP�4weG�y��=���ҁ���e(�.���Z2�hj
�a���ƫ��нKQ�����Ѐ��j,��a3�u-���������Jr�KYG��q�����?�������&|o�N|�#g�^����f� �T��'�-L�S1`5���p�69���C:�x$�������O����i���V���yAuhm>P��	�$ 3mɗ)Z5�h����%���fS�S`⍑�T<�~�)��ߘgz��0ns��c�#�TU�p�R]��& �ӌ>�Nŗ���\a�dSڭm����z �S��yIK�Ԝ�x����t^p���0MF}˻MA4@-���`�P�F��DeR�>�U�h>Z�/����^�u�:���&c�'o~�y�������9�h���n��d0k��!�{.�ߑ|ߥ`� b�u'��#��������h�S�*)���1=Yذ/4����;��C�a7��T��=z��A�ا�����N��a���@R��p��,��CX��㨂}b6˭D���{a�E�a�#�IT�����S�w�
��Ѿ 1M�}��X����˹0�g��_9�NOC�#.��z�y0�B�^B 1�r�Zu���d,.�G=�����֓n�ç���
�d��>�:r�$y��6ꣁ��t��/l9|�G>�<���Z���T*��(
-J�3xG��������Z�d�3ڇt�����Gߘ���?���8�y��wsS��NV��-��s�j�c�L�w���% �L*�{�����!�-K�%t�6�$��ǈ���L�nu	^Lzq���X��nչ@��<yL�(a���H?&��fe��=0����;�q���C�A����yʪ	�jGi��M����y���^.���.6�H`n/X�(��S���p}�W�����(��&bm�����os̓��xDt��.$��\��jW+"���c�������a��	�����8�ّ��xT�3�?W[�M�����3��oz�Wymeڝ�&v|��,��O�/W^A�.B�_���[��+;�TΌɃO�>�+$@0�/Hh���᯳8�Ge����.�O�bg9M�^�����$�밁�������^��#���Q�X��/^���!շ�]�F��ot*�?	@1eې����7;K��Z���;��<#�L5�!f��m�q�����Y�jh�Z��"�<7>�C�T.�b`�@a�l��IUN�Wda�c����24`}�Q�`��D�طK QX���O�M��16�_�+
��̢����&Ro�ﶝ�i5sn�Y�-KB�7��<����ⴎE_��I�'� -��U|y"��AG��^�6�}��:cS����?��ZW��E{�{'E�ܠ����B)��餎�N}���F� ���-a�'2���D�H�T�t�C���x�,TR/M�f�]�2
}A�$�ֿO���7�8gp��s)�v�|�޻!��e'���@I9�Ԥ��֙�iV�>q��(��hW���^�i�������P�>�T���g"-����Ąڥ���Z��X�*:�lQ�TDpT�CR<,9�^������C�e�$�*��F�l���w@ h�sU�dp�c8�>��D�z$ ��<�f�����gx��9B�d�Ѻ�I��]���ob�'��U�
���Q�U�os�Ŏ�b0��򀎂�imz��\�����lh_�1��b�&.gT���"?�6=c�u��
���)�V
�KzǠ��ۆ�&K���%2���d-���0�����^M�^@�x���z�=�F���-��{����"��o$4�t�A���?�4	7\��J�g��ٲ]��qj��י@��Q����P���;DU��.�<�"������vIz��'���U��_�BѶ���	�c(MȚ����Y�	���6����\On�@�n����-��/��yƭJ�)}�&`��jLF�E1eH#���������� �wB�V<Oȟ���F^_�ă�9e�(Ő}��ݝ�x?|�z��J/���R`� =i�@��b����G�^��`'���Y�i)=a�2.}�đ{Z�@�u�EU�.�����i�j_��\�g�L �U�����ɦ؈�\E)@ ��.Vj�n��*�[��t��;�U��TE�0�W�BJ�6�+L�����fPGl��*��L;uP��yɉ�Xn��Q�]�[�E�rŴ{.�O_& 	����+�Sy��j-]s�~N�GSm{�v�SK1���D1��E�J
B�%��~p���1<��!qh@�'*��U9��V�m�����.T|�J1$f����|{D�m�h@��w+�ӯM�ɞ�����ī��鋊�e=1�����/C �m�a��ִ�I��l�@�?ا{AX|�K4չ9�Q$[ev�<�����28sp>	@8�F��~��LYBm���>�ӗJ�y��w�������-���$�5�04hvO�$�b�Qo�uꀆ�/x���(���v3�^�ڌ[�[tiD� ����������R�\cz�-8@�'�{^��"2S����[�e�\��Z�.``���oZ�x��Ձ��e�e���[����S�-9��~�i����t���F�1�FA[}*��o�B�QVt���eJg�)X����T�i�B��l4�E%k�vn�Ĉ1;e��/��b�tN5�_����Ɓ��P����5޿�F�q���������_O\B"�|}��2�	]�;���'�׮&E&%�ǯ
��I�E#�����(�:Y���Ƴ^2F��In�[tp�\D�����e0Y2b��y���:�G������}Ա�?O��Z��g�u�G�j���I��*���1�<�B�W�0��T�K,i:����;�;}�ΖJDp6�^%y >�g�$" m��s%����@S��t]��h��z����̃='ȟ&!�����	��9j3>�JN���Ֆ6B.f��NC����Y9:�꥕X�9�3@��[�l��<eQT^���U�i9�Nu����)琉�h�48��Jt;pJM`1����2�Z<kS��&��bɋ��@������2ng�/l���
h���`![~��o���k�<�Fؕ��1RЇ�Q�k�2*�'?L��kK*d��jt���2n豄���� ]�d6H�����~���!y����I1q:��F݁g.�8U��E�	�����6�Kϡe�*����
&�h�ҁg�F"��$�W�I,a�p�5��h��xw���8V ��H���R*���S���!��\��t,:��rZ�Fz�SK.�-[�0P1��:2���'9Kٔ.��j���9W��O�\���ՓUp�E�\�ʋpղP�@鮎��d��r��ovK��-k�T����=Z MX��,B&IV���}I\|x��_�g
��4�T�Q�yfj�t����遢���l���QN����T<:"?_��0V���\�����ג�5C�����f!���TX�x�$�"�A.�݊�ğ������������>���r����!�9�2����m�E�i9K�~�"��ë��W�k��;)�{4JWN�_�"��HP�*������hV��{�#��>Y��UT���;I���Ź���Hf
(Z��_K'�=� E�^��`"MQ�P���2]M1�_V`#[-�N�e�d!�
%���H\A�f�We�;�`2��D������:v�6��I�p�SՀ��Պ`�{ǣ5����3�,�C�]��w��ԉV7��}N��;�POg5�MPE�pN��:h�#HrJRT���G�*�6?�F��1q�iH�?>kA}��µ#\�W�>�d�����(9�,�.�E;�N_gxGˁ�n�7���tAf���Ƴ���I�Uy�`ѵ��T{���>�/�v��gM;H�t�]bp
��!R���.g�U_���a�����V"�S�N�?c�q*�p9��C<B,�����[ fO-�?�K����X�3� ��������B[�nOܹ��} R�ʞ�
���ӳ�=xSe����r�ZI��S�V��W��`��͑8��]�Y�_׏�ȁ�HR`���p��h���7�*@�L�5�QX�S���0po9fW
0�wW#aT�����u��`����c��(���^����Vs�9�z��u;i� �H؈��H���e]�t��-���Yy;6|(�eh}�4�E�����@J��.�%��.��Evk�(E�d�{ ��V�V&}|��%�	�U�t;F��Qd[\�ln��1�ϖsz��+��$�R���M;��mq�-xdMY[6�8/��H���"[MbC;�u���KA�����x|������\\��O�p�y֗�S^דx�2)i��R%Q����lNz�F��Rye���d�\��y�%_��0��1?5��O�˹���8e��e�P[<l6��7<�%d�ڣ��lv�C��N�$�y�1�i0��p�JO�9e���<�5�@2�*��'T�D���覾�[n.�̤��Gƍ����6~R"u��^��P"�MUwW>�ň��9����o:}�Lwq1:� �H������JԦo
��\���xf��l�$�iՙB��~^H���m�`M�Ak,r�~�^qf���q=|��i����W����>��\�
�U-�1>H�(k�������7s���V$��{�g+��
����\�{�H�P\��O��-u'���C{�ő���ֺ&��i���v'��YL�3@%ґr&:�ʘJTJ�~]�@3C�^� ��/ĶK��t���~���efmh\���w�w	��*�<���&�:Lj/������V�Yg,}�<�Vb4-C:� P0�����A�#�X_�'���	�|H���s�
F��)�NR�HL2��7����*m�Kq8g0�2����W��C���P�i��P����&�����+6����/O{�e�PQ� �rOK*�\�χ�P��~��0ԟ"ojT�'s�.f��nϡ <v�8�/{R)f塚`�T�����uXV}b6��;��,��dw0�Š�N`J*��U.#�6�o��(@#�ա
�b�2��F�|^�7��(�ل�_��%����t��J�Kdww��і}�ޓ�UY:ܝ��� ��}�Y&ߥRp���ޢ�o`�ª��P:LZ���]I��t�	�.�(���_��)z��"�p ���p���"�A#8�Ue컶'8K2UE�B��L�1ԃ�n��6�0e֯=T;C[0�CG03��D��d�D����i�;��Ցl8����o��Pv��L:5ppL+SK������n��2�P�����3�L(6� ��L�v谍i`ө�']�X����%��x�H�|�F5�>��Nd<��#��l����)�eh��t[v*4���q:<e�JpF�4�Ek���{����~{�x��Q����z��"e�dp�\힟�Zj���^r���!�V����e|�>x%����ӱ��}�Pv�P�P�2�V�Y$B�5]50 ��m��zR��>'��_˥� �=�xi������\��Yb
�ا�R=RK��T=������y� �A�\f���W�b�!o��V���2����ŀ��|*�M?��B�TY&���]��ޅ�}�Ay��X�Q�C�c�����s6-k��ϲ1h���wTc�;���fVw}��W�>�a�Ss��1�S.P�
ɣ6�???V2ނ�����s���#��6Lf�fu
+l6�Ɵ~�� ��T��X~��O����m)-L��M�<�=�!&�@�D����_H�v�?�8)%��L-������J�^[us�Н�l�7)K�U��ڬt,�Z2��pdR09�K��~$�א�`=zX��9N)�w"�>&��q���$��]-`�s֪��Q���x(<�Q�z �V҅�$*go�E-��D�(�e��R3��&R4�^�r�)E�w	aƁ��y<���YY�5۟���{��u���+�d��Dhu>`�X����^І&��gT%a�GaikQuP�,�?�oH�%�j7aL~t]ew3��NJ���=1�	�|�曌�����,�5��]~�-[�E�%���Lf��g��e�Ɉf�T��ޘ���K��G�%(QL~F�"E$Y�Q��^�B�_x�X�� .�V�Цy\A�T����e/�/�?n��'��&�-.��Е�ƔZ��i	S�D2� gJ6be�sÄ�:�a2x�,v&*8���b�zT����m���i��)��þ5' �}��T�����\�q���	c8�s�k� Gt�����6����RS<?�NT]��1��lG�j�����~G��q������S�jR�CfT���y�,�������D�Ng'��B�L���H��1�\�P��J�^Y���^{�CY���Jy1�?z߅����Ω��h/����m
�8|�V��c���irg�-�:�i9)�����:�A5�C�C��n/J�n�MVY�I"������}�:���"�-ٿ`��>��񨵽�%�ؒ!��'�`�P˃}��i`x��A7��w�nB�H�
�Ƨ-���_͌A��r,��G��ׁƈ�I����;RnȨ��w $��v�5پ)��ߤ�X��>Fi%�|��5R�	-d�u��������	A�'Mk\��)����K�c� ��YX�g��n3h�%%:���c�/G�ĕ��0�͎pmf3K�G�m��r���Pe�cv�|˽���+�rp�5�v6t/�5Z<���QƩ�&�.��ڊ�����1����1���\�4���v��Jf��oz�@�G#7��&2����+�֩*	�~�A��.=ƐC��+C��s�Yh����0e�§���ǔ��U�э�{�
"̀��w�\��h��`:�J|fs�ƙ�I�"��8�N^O0Q��U���F�4(�(ހ�kyXvR{7/hg��#^�>f��]��(H�)�b	�6���������Jꉷ�w�-|oLTZ��c���q}ZUR2��_�;ta�j6�?+e�0W�N'61���K�]�LX�j�wh�*	�)��󞌉�t�.����r<�2�N���������)w�/Ѷ8P��K\�����Wj�|}�Y���{Y�I)4��:~ᮊNݹ�+�����]�=�0C�0%>�:5ew�P��XW\:	#�kh%>�Z�3�z��i�i����BiU6|��� ��X������d��k�����YP���=�5"F��I�ø|���s��~`0b���){s����J�A��#�V��g$���_�-��U�^�)�Tճ�U���4�@dUUiI���I�8�\�K���H_�d��7ɥs0|�8~��*y���]al{hfmw}ߦ\-?�V=�d�C��o��h��&}��&jr�KzyG�x�P�_X�[Y(�m�6�&��&KEd���O-88����1��pX�=V<w�����iX��$�1�O=Db_�h�
�<�m���s-�Ε�6�޲B��H���
��Lt��5�@&@>ꖣ���u���C���BKDi��2�#���,�(�:CE��<ݏk���~͝g�|��u�r�/meT�Ge�h3��8���f���.����>�r�Ď�*�ؽoZs���cː��i���� ��t���l�O&p�#����iX�<����WR�y�V�N/���C�Og"Ϲl�!U7���^�%��Пmj$�I�+i�U�麚ԧнE���c\���T��ŀW�k��z� ��ˊh��£FI]��+X��X6fϩ��)z��|�q3ݘ5�L��r>㮽���+���B�m�g�v��J�,86�$���w:y�`��mih���7	�y+0yY�V��M��S�2�*B�����佉���|@�[���iܸ ����D��q�d�F4X';Ѫ�4w �[Rʖ�:���/ˠ';������C�j�e������NC�`~�_+���EpAW�4�0���[�΀����!W���E���GYfؼ���d��P2�H�����ץ�Kp`Bq�PgY�	d��@@u)l6!V��	��������sy'4ׯ�z�4
��8NQ�l��l�qYXa������U����)�/M�2t����k��V�}3n�&�U^��G\R��#�LP�.��	��\��v�V_���BL1ק%'I�b���ͮx�������:Z=X��x���*s߸a�4�m�0�fy���Gv�d
�$�'[DH2M�����|nu+��L��w����!��Q�(IHS�pT*2�j��d�{��pT5�^	ȩOgk��ٗרl�ާA#�e�̡��HL��{�b�]�H'ߐ(B��t#H�n�&	�S;I�z���%Ǡ,#ӊ��񈃂�a��W���!�0�8�<�> <��{���s�����+[�#R(n�U�eN�Xf�/֤�s�b�3q���)��KE�T�-y`7���L�1�[bJ/�x��	��zp餻-9�L&k[)�H� ��Su��{6A��C�ٌ�	
�i%g��ekPp��`z�F�_Y�fY|�#?1�k����.�q�G��g���r��ż�5*A�`����@]?^�Q�FY��H���WeG{�v�v,����"�}�m���d��e
׏�#6��@���W/�e�+��QL�!�Hg�ڑ���AO4:��`b]O@ฐ���>���w;�QA]�v\�Vn醟F�-·A4�DF*�MЦrŐpK[^ĺ�[�|�2i�>@	�k5��m����kKO��J�;�V��+�N�h�_�A@q���&�p�c38D����!�{���F���	3�CJ�yD��Yi0����VA &�ގ�����V�L_�U�]��=}�,���'��ӺQ���A�Դ�r�IY���M1n����$�"�/�[%^�j	���?��)&1�5��1c���jT$}�W�\H?�t������h;5�%W��"oBɜ��?t:��P��x��0dl�ç���H-e���Uu%��Q�@&�)�Cz���l�ˀ�\��5=�^s9�= y�����zR��Ղ�G!�/L3u�^����'�4�	+[/������t�ZP
'��`���t�-P]�ڃ����$��c
s�n�#N|�R����ZY�����<����P����1��Z&��%n��uY�A�C�fT9�!b��֬�.b���P�!u�����f ���@?o>w�S�Zyt����Di�R_��Zm��S�[Diϝ��u+[Ȓ�Hޫ���d.	؜�yi��P�^{a�~J��>�� 6J^i٣ˉ�$���ޮc{��4����N�V�4UZc%k��@o�și��%��
��T�S����۞
�4Z�*�qf��C���łs�+˖7��V�c��R�g��M��Z��4��^r	H��WA���a���8%�0��'8�ˡ�Y���K��J����a٘$���y\v.��e�7��;~{�H�%�(^Ejc��y�Hמn�{,���mߡ[��a�ƻ:كv� WZ��j�b�o1�Q5JQ�lM=&�ޝl��,���:@��h����oO������±~�Fg�FM���=R<�Xr���[?˒��2�U�����مWY�`�u,XBRA:�{�{�!��%�!'��� ^mNK9���o>̓C��bY+�|
�ɀ���[ܠ}����1Pϥ$U�B�2��V~րf`�)�J4TU&�P�hb���h���ś�_�_�K�#�b8��n����D�#������ƲEN��'�x|�m��3/���N8?[~O��kz��/�5.ͦ����1&ڶ���.7���Q@/��qe6��|�Q�p��Ͽk.o%@��*�6��l���S˅͸ݝ�-�"��=XhtKl ���C�YPH���������z�I�y[t�Ƒ	�v	�ۘ$��B�n��qB�I����<!��笏X��c\v4��P׀:+q5_j����e���hǀ\�>�kX��{�fO"�о�˜�O`��;.�K��Q@괟🠴��Hi�_�}�&��5�N�����1����3 �����S�\��M�
��񥥪���zP�2���m�|��D����^�ǃNT�6\5�<E)�����`�x.�Ǣ��_��S����}�	LO����7�k�3˾�tz�x[�&��پ�!���pYmR��q�Fm� 029��� �/3����QI�����ZqZ���5j�����bƪ����/�b�O�4Y�zJ�����Л�ش �8���Ha���O�8�׏@�z*7
��?�o<iM��j����Əq(��lﵴ������M7m�,�\1=Yu��O��u�a�ݕQ������;�/N���p�3��E�y����[@�^�C��U�H� �2�f:�)3F���$�5��@+͕d��N@e���ި���֥���L`��n���R�\�/(�<����y�&vE��?6X�Q۩z��xA�p�/!c��s)v�3q}�1[^�o!��F�ÚY
#�5�gb׀�s��3�M�����+_��c0S�:��%��Yx8�y�t�^OGx�5�����zHBX�=zH*��>�cVMb��z4ֆI�\M� '��՞����cy7fL(�O��2��;42��-�o��C�������1$c�9�ٲ,�!}�f`�P��}�co`k��)��D|�ltd����v̾��c߇)�'���+��RF��v"҂��!��4P�:"p�޽�LQ�'�hr��v󣃦U����:Xk��'�

���?�4K�}�9M)L&�D.�����$�n�AZ4��-�z�v�gxf�4�2$S�R�O�	�S=�5�	��ȴ�_�����R�O Ljk����N)xˬ>���Z�V�Z;�):�1�E\�x6k������I��t^��C��k\i�-V锚�a5h¾'�;H���4Z��+~4[k3G��`���L�2n4h^�J�^�6	��
�dA� 5Е�joC�@�0j^(��V��2�;��D���	"�
X�(pro��k*?�"���~FaH�R���XE�*g�{"�J�~���װJn�O�&ĂoL������:�������L�oe���y���T����Ͱn׫��W��+��X��g��
3�	�ų�������&6~jC��Mwc���G���Is��۫3ie4�>������u��pn�^�%��D�r�#����*�T�-r�G�i����I�i���*�q�J5 �v"������N]Б�e���w$H?��T�,����>)О��F�\��Ѱ�4&s�꿟��*Je;+��6��TT�
�[Z��GR�I���_���s���0�|�eU!���w��l����C�Ds#ݏ��֦MT�%V0����6�ԫ�wD]yV���bǊ�����l���[�tJ�vź��G�;v�B��*nu&�Cѵ�$(�.!�#����g�Ѯ���y�T7�5eLwl��sWq���w6u�dԗ�R���8����oӂC�������c�������=�+������R�&��x�1$�ÿ��uMSXT%ߙ�R�7���Ҙ��>3�PBB��!���(����i�K:�q@�0ki��T�<׷�jWv��i�o�Z�9@dL4fJ%t�ܼU�x<�5K"�ߝv����<�"W%�y��:[�q�7��"�kfH,�Z�@B"h���a���M�s;d}�q����a d�c&�D��d�f� {H���U�#6>����$���j"���k�-Ȟ��Iz�c�h�ce�H���/}�i{���Ӡi��?��H�.���GdK����0��t�@�I���Fj��	@��{^�*B�7�	>M���6r�D���^�x-��kU��r�4�1�鏮t�@�ͻ>�ya�f��Ϛ,;f�9�d��C�<ja��=��t�$�E�cE>RL�Ձ=˩0�H���4@�;�j�}���uM�nS�v��!��5�$35�S�r+�&���S3�R��vI�c7�cC�Q�Н�E�y/�ϰ�$��%�V/� �j�;W+��n��iy�]�HД��b����,�:�,����u��T,=���Bp˄<٭����7�A�$q0�9ȯPw���d5?�h�/�a�)��p�-��ء�㤫1����
\.9=J�Q �HTՄc���߲�ѷ�t[�yB� 0�o���	(W*�^.lW2��U��ϳOI� ��{o�; �JŸhO���X��=c' �%(�?��0�ʵ7)$o�����Lz�b$�,���C����E��:�8�P/�6~�+t�� RӃa,\mp���h��*�ǲˏe�&�X��W�C�h-&]{���*�����%���ا����1��!b\�64�������Z�3؁�xpXqk��u�V�_֥&��#��j7�v��w0�Lw�0��[G�g���_Rtei|>���S"�ʆ���fU[N�ee��_L<L�U�@��Eм~����ӟ���	�b��Kw���v���Q蚫��4��}HeGE��%sGT1�L�3��] ��`Y�f�ol:��{3bg� �	�����b�����-n7AT�6��8��S����ƌ�OQ:�	�[sm:��7ǽ�'�r��)��!��ZzI�i
gc�ç�i�pX���_a�dO�, (�Ւ	��#�y}�6�]��LYOW�هd��N��F�ZU�V�	zNN���!#AĨ%$I�t�<C38vI�����b@���,���|���sW>p�����ѣ
i���%�oe������J|�ԟ�#j{�>���C7�iA8%�����F��n�#Gox~�{*_����-#%������2��>u�2>V�Mk�{�U��!����ը3��?��
����D�(�!���uռ�lä³�{y�I��r�ό?"����M�k�$�&���5�������J�IY��##�v�6�I:��	��RH�	T戻���l=ʅ+����_�Dml�1��"?&+��=�N��o�E�d�����`�Xθ��,��[/fwy�,�1Lm1V�Q�� %x�*�<1��x�g���6������!�K��dOy�O?y!ֶ��xs��[���笆�gR�S��;  �2Ŵ-E���f��f��2�G��0�]�6_j�-�����o��g?����˃-�'��U�:�!>�_�Uu�馍v�`;P'}fq1PP�+?��(���7zGo�-��ź��.ۈ.g,D2��SY���C����0�W�7cl3���	��Z�$E���?�꼫�6
R'��=��Em����1��s#�}SX��b��==c"Aڮ�E`���ޮA�(q����g��hǔ��<B� x�$����'=.>R'���a�?
ŀ��~�1�60��nco��j�&�-�7��4�I+��)}<}u��jQ�b]��|z��)���6�C!J0ʞ���9�iɮ..C9T�7�ce�t�R��z��mi2�-��:ʜ���"*BHųc�o�>ˠ���-�\g��)�ya�fZ(�������a��V�	���Tȵ���1���N����&9��2w�澏f�)jo��:���]�2����=�%<_��R�#���h\���EO�����K��p�F�����U�'{u �
5u���z�2ܖ�؄�:f���[hw�#P��ѽ�L�_��f2k�U�GD����D�P����>a <~�CHcHW�y��E�[� D���Lm�P���Lv�mA�l��i�����:#�V���,��%s7����R]ȅ��E��A^H�Xe���I�3dէ:q{!r4���`���6����n;[I�'P�Ɂ,x5��](��9�eJ �O1S3��
xq�?����)KՋ��l.��Â-�)�Ij��΢�޹y�Ə:b�w�q�GO��3�Kn췛�`v��7������L�MQ�e��^�[`�����a�ș|����͢��C�\��z\ui�@z�P�-{�eE�R8�����|&u��)^�a�-�_Έl;}�A�M3���"ɑP��<�t���$,e�ޝ�F�"XsD`���I������Nx���qPR�|2e����� 44�i%%��xO<1�Ĵ�c�>�T�>�ˈs�F�X8�-t�Q��@��<����E�n��B�ϱ���#v}	 x���8�?����(u���Qͦ!�>����ѧL�=�=4.��:��K�\��zԂ��Ă��FP�mvNHlhn�?0���hs����Z�/A�?W��G��p��<ޓ�vemj��ܿQ<�I䷿�G��٠&�W]2��?��җ쁵j�WM�j]V�m�m�s�aVh�]G�x����z묑��R���0E~�nK8�̅��'�3�]���*\S@���d�9	 On~M��f�r�5� �>[ޜ�-�`��|_c[U$2���K�(r��j�'s���3���S��_�(�΢�������(�ٜ����=\��K*�-��m'7�r(G�d��-��暶k.5�V�~:�����V��,���R�؉�����R�8��K~�4������h��\��-EpDDw�əD;��	�	��X ԥ������؀��<�_����w����S_AѠ.�ytq:������RGL��a=���⮓o�N߹A�S��ҭ����#�G6nS�>rM������h��Kb.�Z����k�DoFՊr�&���f[c#(����5�M�zŌ������$A�(����3܉�����i�ݍ����W��r�+Zc�|�^�[N �ڸ��{�^6m7p�O��sSᠠ�z����Ș�c��Pv)6d'�,Ѯ� �i�O1���߀S�kK�$�k��Kr��>,dVL88����[v�������ox�zDeTˍ�r��#���pjI�L\L�r?�2����3��;�W@+���k��)��ۜ�U ܦ�|��RE��oMẍ́�0����U?:{�";�14�{�6E��T�`� �i�Z�Q����v7��%�c��{���q��4+�v�[�"�Lv/�~�u�uZ��3w�%�7S��@� X4�_�o�Fc1�����Y[W�5����y����:�|>ƭM6'@�`H"�x�U7�iT~����NX�O6����`���^	rP�J����k��� ��;�����"�\�����g� �b�4�=u����L��T���XЄ�"����Vג/킒�( W��^("Q�tCL�sEHT�Sf+�"�Qqp���4��-I��U��t�LH���HA�o�0,�ݏS����|Y��ݻk�r��Jn
�>$e?��h�;-"��p��+��;�VF�.��W�jo��-9�@��oP��5��/��{`�z'j��Ė)�q����ۚO�_Ϲ&��~��ٗ��Es
����l�Ah���Ι���b�t�E�,�El������X`�1mB���<ԬG�j̼�;�&`��>�]�����ѕ.�MwDZ�G���e���\�ȶ�n��=�jZ��Wk6��E���;DNH��Z,t&��6v�8����KN;������b�|����XH����n�H�P2M��&�؞5����
���|B�*{5\N�}4��BE�haW�%k<ߦ>���3(�XS����}�K�[K�ΖK�A�2r�c��}��
�_-0���0��hs�b)�my���9���<��`��㺮#�ㅉ����!�ER��1�J&��X�<'��y�\����
f�aR�n�F<|�a����"h�)q�RZ�Z�DF??)ZN�b��ڳ�b���8m�্��<�>�N����(re�ի�$�Y¨�*6���������&�N/����+pf���)�.�J��	��r@o_��N���:�hg��1�c6��Ss�ދ$����@vA���[��b&O
a��;�|�r/�NN*ҁ�y-@�n6Gv1�)��K2��q�)K1�t@W����k�$x�;���H+�����Ա�o��Z�]�D{ݚN.�n�5K�W�_�5���|�6v2�m1��/�<s]Ô���j蕺i�g���p���?��⸩����N�����ۙo���V����+\�}ƀ�Ko�i�O�����. I~��Vwۿ�ԍ�+��Åg\�e,d��`�]HX9�Y̡R���&��})��h �*��<���/�ڣ���@�-��\@���R	��`�L��َg�zI.Cpya��I�m`F)RN_%���/�����3�H3��1��A�?f	��<�0�†�`�F��9�Er^5�7�u�1�����ۆ4��=.1M�j>k�9��S+F���a ���R�|o�?���T�v6^��h�0/c�T~T{j���{_�w�sa�'?��n�D�w�r2�I&��B/�\ā���)��/�L�:�@(�����x���S�x@\�g�m9Y��isD��{�nMo�[�0�򚡺R���EP��Q��3��J;���ΓfM��V�{��i��8����,���}�m;Q��i��1���2LJ��9��A���}k�A�kDJ,f�,S��TqyWY��#z��2�8+Ԭ��k���C ��X@t�!z�p\2��ŘPѽ�I-�ɢW������$$���{�~� �?��Uaj	ܠE,)+��i�/]_��� `s?u����,K��n/>��r�g(��q$�� ن�R��hdP����>}'t�^�^ �a�y�SA�^8���y�������^�*s��W��q���h�Zl,Y�����!hѕ��:��׍Һf�-v�X�*��4*bZj����o9*�<��-�>^��Ą�B�|��Y��&�-F���_�: Q��{"�FY
�=���Gc����.0�Z�3�i
Q ڑ�7�_�C}��XWK*PD�A�R�H,�`���ha�r�1��6���U�iD� B1�鸃�h�C�fRU��!�=���� M�cdQ�at�l�V-L������8rW30pV�+�}���v���-�
ö�qMB��5*� ե���yFD�	7m���U�ğ�ڝ6�'^��6��}�D��~�)v�]��jI*�\��ҁ=�xY�Y����1����+4������������U}t��N��Y�7Q��Vq�� }��G�8��j4�"��O��-��N�;��S�YA4<� �q$ʙEl?��o>��h�0T&�fK?��ij�b͕(b���%I��RXn�lq������n�P�{d^�ԫ��ܘ,pdޱ�ʿ�7VON���a2К^�ue/�t}%P�cz�إ��rZ����IN�j�D#&P�xن )��������L��z�%��C-6��B؂�y�z%�J�cU���Mm����	g�6���Ej�5(a������1��V�����~R�l5�d,��m؈	���C���K���y��=8K>9�A�.����	�B��c3B���i�k���{����?Gq�5)����Zd�D�(y.Ns;�tK|�"��|��O�'	��3*�]8
�.����|�����_�˕�����b�R?�)d��856��*���֖�-3%U#*�.u�$�ɛ����u[�S��SmBE���!Y%��
ܥ�3"����9��I�'�0ϙ�����nҦQ�*���]����R��&? �����A�1�Mb�T
3n3K�EB=���U	$w:?7%*<���0�hҗw�ʿ���D�u.jl�*|���
��j�{����`Z������I*h���l���81a�S�v�D���k�N<=Eu�)1�?z]bPVx{X5��`�
�S��bPFz�۴	P��.\��D.�������5� Ν�y��ڄ$��h��?Hv�p����IYߗ
�e�� �&��Zcv���b���z8Y�����p[�
m���x
�K�1Dr0[x��k�aRH	Z}j����V.�)Y[hp�����ޞTI[ܫ� �J������mɔ�5ԡ �]�����b����y$����N?����A	�ڽ1��4#�Uٸ�z�mh��=�>�0W��b[��D���0�B���������zL �~>��a})C,W� XB%u��)�r�Y�f��a�mr&)x{X�+l�Aj������y��s
�%{�nD��kŗ����� �4L�c�-F�Sm0����)M��
��Y�	�?�τ�^ɍ�՛׾�����\A.5�j��خ��}?�.���ʔ)�	vFW|��L>����x+X[�l��p���vF��kJ�
��*أ<������sq0|�&o��n1��ZH*�rG�D�u���c�����	�Z&܊��O�V�~���p?�x�U�GuFQ/ӧ���i��m�|���z<??��j⧦�VzO����8�Ұ�Qe��mD�N���x��9g)�^sf/��~![�I�u|�d]���R�4�N�$�4�%�I�Y�Y�%"�GD��S��L�����'gf�X���l���H�-U̅�L�ڣ�JO�ʒ"���������#�#v`����$dN[�ٿ
��V����qe�K�Eh�cQ��<k�xOR��4 ��	��Rm�^�=,K�R��(��xr.�$	1�e�W.x��<U>v�7� t�5��f���9�OT��i�z�l�;�'��O?�w���%F$�@H�rY'���cAw&W3|����#�V�{��.m��7(�n���P�uG�^/o�����@fPp^''c<z���$�Ɵ64Q"�ϛ�C�e�M�f:�s�U���ay�h�����g��ab:�K�!l�iI���8ZW���"�{޴f��s?�EP�I�cܓ�󉗌<Lv��w�wپ˽2<T�T�Zk����R��[{	�RP��X� �s^ی#�+I��m�^ ~��������㬂��S9�Rx���X ������VZD-/�|C���$�s�~B��1��hw��̽o�%HmM�s?�)mk��1|r��m���Tپ�k�Pr�� �,��r'uX��B�	E�M�98W6C�Inf�
��'�1���bd����02q�^b��l�o��F)���ˌ����j�����p{�u���r|`�Ҁ��ak��JN>���t��`�VӶ6F�Lpw����eˠ��<��M!�<���t��1�^@��@�9�ˎ(��JE�Z�}�
�cSѴ��������z�)AiX/���؜����SE� ���1b���[R�z�b,���|�թWh(���7#t#%8e�w�t��E���ނB`ڭ���z�6����ai��M>>DN�s�]	$�9�Y�������z�M�z������ܲ@����r!�U�A�n֍�����r��f/x�u��%Q'uY�(�>o�x��{E�tY���rt��=5��v�\���7�|�.vx�#�(�_g߮$ &8�"6^��=�
���Q���|���=��O�oE�I!H�����	ل�B��b�'��to�{��'ἇ�Xh�y� �BC��)\&u�W�?y����[ #�Ht���GF���8�9܈�nplԪ,��Z��W�T���I�]�
n�_ӇK��9>�fϻ�o�D'������~�h�Y��dR>��jq���os��&��7��b7�y���"M?����Y=0-{w� ]@?]la����x�;�[��-F[֮�5 )NP������%7�B�Y��0]@$x�KX���Q�y���Ԍ�۱�����'B�K����4�����'b�Z��FB6&9��S+�S��TP8 fe��l%5Q|����,[V���'�G�+���}F��{�y�Cs֍���]j�%���<�Q��}�^�����S9�C��z@Gc�5~�$�~W<1�֖�����ZїqU���:��FJM��g&��G1*C�]�OF�>@@j"y���`��f�:?ӻFJ�6Fd(�X�Fw�O��r �~�<�??�&|�F�(]�^�G �'�+� �s�9��$	�k(���M��=_1X���73H�cLM�c��P>]�4��:3:�r1�`葪�B^�]^&�l�7C|�g�w��u�ڔYW�a�;�ܙ7H_�����n6�DΧ��)�ҍ����n ��]t)�&�еr�*C&B��E��}�<1��u}����ۦ+-M7X5��;}�,j���3V�U닦�c�T���b��t�qLu�eX.�:3tW.�j�	w�}1 ���
�=_l�Lj�^���5�2S�{^̪�O\0�N�&d�r�Y��=�OR����x+����K�8��F�J�,��]Z�6����)�LKs����3(�����'��>^��+6��Ƹ
寎ʑ�����ԏM��C���M��O�rP`�r4�� ��T�5�l��Q��TTR��*���:3���?Ns��q��:�H_����$s�����/�Jӂ�-�p-|_<V����'1��wy�c���,Σ���@-P��g�Ϩ��v���D�^�J�EcB9�f�`�.B+��G���	E���,�5N�ҧ;Sh'�m�~�����u��%{�WQ�Sem\�flC[���VO�u�K�&	�ۥ��t
o��'1�K�<}v��58=��s`>/)����tjN�Y8��$ƭ�N�l�G���5���3�t�k�6�,?�3K�E������NSz���PfwW�MWX"U��Hî��,�8%C&�[L���{�k��;�P�_��}���#}�Givn����b~$2��/���/���b���`u�ʏ�أ�QP���������u��f�r�k9�}��#JD�3���u�F�9��-� � Gy��ߖ��B����9�O���$��k���-K�3�fۀJ<�є�rm��X�����~���Tb���]��gW�`�[HCƩ�?�	P��|l��
�S�>(�I��E�����#��&��O���&��M����r��k����AD�B�΄�[	AZ��e3�܃����zk��K�t�f���;z0�A�_%C���!7�k����T?-*A
��u���.e�_���m��id����,N<�ӧ�y�6
8��g॒�h(45m�>T��74^����N�������A�U�w (�(��Gpy+Ɯ���/q�-�.sQ����_a7CBN����� e9 �H����waR�1�y�kx�|������d��$�F�Y~��Fb�OH�����!#���;|m�?@"�C�$�c��.=E�习�{q���g�9��_'�.�_$���]���#�IS)nFw�Ƿ��m���=�0+������v2��-Q|�����ʠj�/ __+<F�΃>a��9&2��LR ��PX���s����hپxf�\�����n�wv�p�jN��B�U�Ju�;7�$�]��.�Ҁ/K��� m�*�]p݌Z~�6Y6��J�Z�ш�ǑsK�i�������/	@WNZ���a�"-ȓU���U2�L�B�UvP�����,�"ye��u^|���&�f�	��~j����5Ia� Z�憞�ը%��0�鸕J�E�v�g𣒟��u�d��A�qi�"H�oW�<*����A�K�M���1ɼ�`���@;mx��Q?��=��#�uw�q�9g8p"P����㰣���!����\dK��KV�b��G��Cx��99!琜J�KnL.�]�Jf��#0�R[w�R��������і��9l��󬏹�"�r�ʄ�l�b��4��Br/�6f�dy����~�B��M�P�^5�J��eĖ��P�g����{x��Ȟz���f��,�J��Q�IED�p־P�sf/��� ��j��T�2�η|�*���Z��LU�y(���[��Y�8�wc@N��H"�(c�"Ċx�I��ٌI�f��!�hk��ӻdgЏ$ݪL�E%h�ȩ���k�-~ڏ58�l�&|���/�7�V��W�j ]��.���4׫��[@:�Sш�������?�b��D�Wl3vy����s<�#��Z����
����y�Q���f/�Q����+g&]���+��/[<���.�ae�*��rA����F���`?<�J{�<48�	0sż�q���PdE&�)EXfi6� g�?S4(�t��5��7E�62Բ�uD�JW��N�\�QG\a�� w�	a�$z�W�����P��}�B����P��_sSe�oK
u�U���گ�'�;��:�����m�*��$� ��kh�fU��c�>{�Lz��)˷Й���]9��h���&����ɾ����Z�]a|�4��
�,�-玒̆,%���D��o�CK�u72Z�D#(�ψ�rSQi���\}�7���p9
�.9�i�(�Dt�f�E�G
��ЀCu%*�4���eb#����p�H 2f_������,-6��d�K��-�=�ΰbKv�5i���'E���&��@�)��[J�Y�w;��x�y���E����j���r��k/�� �
���Ƞ���k�@�ͽ@��V�ƃ'^\K�r��-��N68Ep�j`TF敷K��K-yi��B�еcrM̱d��җ�C��T�:�	�5#,��UL�\��=GyGDM��-a�����'P�:�R�Bxb�Ws���N��N3T2��H��Y)��=��I������ ��R�,@O�PS�޼���ECbJ/�n��A���t�o�ƌʿ��)�$\�&)�Ďf �3�0y��/!"����c�g��w6��PVd���,LENWǾh��Q��d��e%3XZ�����TT^@,�p��J��ȼX�h����T/��
M1���J?H�;i�<uMl�bq2�ϝ��jR�h�Tk:��[sU��<��8h�ľ<Pl��2§�r��;3.;��9�*{a�@���Qk��J�(���οm�l?�crP��2�W�O:?!CZ��OU��:������w�̔'��dcҀ��}����	��N�l��'1I��" �ɏ+D�c-*ox�_GdM%���+]� �{�6x!F�ncBr���A	μ�zϼ^*ol0�
2��D#`0����~�� ��T��F�4��	�-~���Rϲ�.js�$�ͬ����Aw�~?W�
�]V�>!E���4�H(n��k(�;���I�}>��'���}�B}���������|��X��q���}��c�ۧ�.�2��g*
8V4tG��ew��aV�#��l��d�𛑤�����)�S��r@�P�Y����M��(g�P���\��G<�=��)��"��'xPT�a��tl������p�+F�F)����Y�z&Sho�]��1�[q� à��N�7�n�U�d ��*��;������{˃1z-dɫ�ܻ��/�9��!�y�����1T����T���t��;��H��N/��d?��J��r'�h��\(wyͽ&p��M[h��!�ӻ�g��=�q�}=h�GE5��e��Hx���g�>D�3?�f�< \�8y��$���Crc�A)1��t�f�׈�7>�u�����s��	s�� O2�mg��a�}���q7�t��}3�e/��ܓ�2�\�Y�p_�eL& 5����w����XT^�%@8�x?n�y2�W��gX	��Q}��[�6�!�iL��M����n^�2���.Q��)��K�C!���%� ʍ�)���V��YS����?�Σ��Ű�3�in�˅O��&��zPZ1Ů�4�_)��zC~'9���Vq-�o�wW�ҹPDʯ5�W��&S��-�L4q
9Nj�G1s�"\��>~c^Oi
�pdSW�:��;�Wͫ�~�ƚ��܎���R!e��b��̓b9��{�'�d��J"2�����d���z0�O��q6���т�� 
�ɰVg1�NSx�@2���"�#�b�|	i�OQ/�e�Z$Xs~�A��!1D�K�	�����ؕ�P�s�<��8��wƜz�iJڢ�·dq��]����P�<?f9|}��H�ܭ)R���U ��������:�S�9���
�K�R�$�7�ݳ@Ȗ+��������MA��צՕ���lPt�^p`=��r����ߥ�����?Ju�os�˵˞-{4��4g7��aEP<�bu�6�߼/� //�P	��w���pi��}�&,�>��U��u����l+�,T�_����ݘ�]6Q�?>���E��yJg�B�y..#w�G���<�U���aH����J��P�^��n��	h��o��ڶB.(��;%^I ɅЙ�^�G�� ���M�\����zǞ.@k���Qam�g1��G ��TME'xpU�ʆ1<�s.��m�/a�\Ӿ_uLvo�=�9�&����Cշ']#�`����G..���yw�"�}0�9����f$���jQ�<f���s���c6rl#78(��>xރ�,l��m�e�Xg��"����#>��V�����S6q0����Ԩ�'�"�&/���~>�ڳ���؋���eR�ⅈ�
���^�����I�ϥ�Þ1.(�{)�:�]ft�F�óت����9����� �5�"���b �o���V�^��`��J%a�[�T|��������d�E��]��Mg��& &��-�+9���9��;�U�����)#[/w{�-/�6e��[�nch�]ו�s+\�x��������];8�WD�0���ö�YG	S�EAl�%�3@��EI��O��Z�~h�ٍV��0*��@04 u���VJM���f[׌�|h�*ERs�<�]:��]x�v4p�@�<��ϸ���p�t�r�w�͜��ݱD�ED��x,\�����5��M�g�n�]�Q�)j�L�^�z郿���\�@�$j��Z�����U�v��`N�-��H|~����3p������	���C���"{o�O���~�c	��Q�� �A�!B�I�;�԰�{tU�&���2ҝ�*�;煄{�0/Ѵ�-�5��)DXgM�>��)�FSaQƀt�ma(0P��/�r��Y�~�M��HF�Ɲ�8��(X�ҾJ����7�P/؉�c}ײ�w�ЍP&�����"+�X�@�{�8��,N렺�)�9��H����>`LLT����/���퍋�g��/�q��=�&��EM��/=|��8-���3r��?���X�oI������6�� U���W���w�~w"�����2���!�y�+�S�%����P����^A���������	�۹�W ���ܪ�d�<��͠�<J��!��l}�\��������ac� ���%���6#4@g� �l~�
�1:(�#���	B����%���uT@�]��6RC�_4F���e$<�e��,>�j���d���Su�]�
퀣~[�NI����X��i��J�����#�Pu�ЊV���<F����3.{�&N���NJ�fk"g� ���~1���C�@-���k�2P%�c����̳�n8/�J��ot�f�X���;�>�M���0X�<��7v%�`$�I:����ː�-`Z� ����L�X[iw1�4��L�E�<cK���������c\��j/��⦕�t�҆L�Q��f��\ ��0*����<6�b�4W�uܿ[� �-�4������Ec��*�4dL4�W��6��;��6���;�n��l���|Ԩ�<����Xu�ȏ+�w�F�z-&�
ev�f���/�i�XHP��)fr��P$\�}7ih�i�s�G�g�>fZ�hގWH�ڈ՗�Q><5A�N�����Bh}�������d�i�!�%s��{�#�^���������;�ǅB�ȓ����Qڵ��`�JE���]�����Z*m��?[����r2�n�h�Ҽ*��Q�Q��v��;Q>6݊b��}�!�f3��<Td&]�a���w�:6��X��E�N���[*�r|C
v��q��>�Eߊ�	^����S�:J�E�����g��Z�����XL������J�␁�\2�^o+
�-+�����ksѪ�;y2���^~|E�������S%��qe�����{��C������X��!����2�(h�\N=$;"�fw1�߂r�s�+��\�U?��'��ԇC�xXuA�����9�����Dk���:��;�|�!�?d!�}y����+;���1���$uG��`JE2�3�:�N�b�q�Ҵ.f��k�v�[fz � -ϗ+��t�x��@<�ޕt[�����\��"Oǥ��e.�]��f�񇫖���HWjh�j�z���77%ݒ,7ĠI1S=��94"�h���ҥڻ�Ku��PIR�Y��PRs\o� ��c���p���+��q��'�V�<L�E�$0}[I�3_=��U�z�q��N�3�m�[|���Bi]v��Xb�v��}QX���H�Rm�50Em�(���U]RB�`[U�p����g��g1t��;��D<�=ʸkԤg�ƱH��dA{��&�7"����y�����͂UX��n}L�yPrw�Ʉ�ߴ�P���1�Mlv!C
��|�}O�Yn�oRO@���6B*�zƄ�=5+Om�o�O���Ŀ�6x�pԀ��@r%st������¬�?ީ�q&@���Ah鎘=+$�_��lp��4-���P���
���i~e��$(�1����-B兲�h��i�.�*R���k�($ՐAǵ��6�z��ߝ�#5�<Mg�Sگ��2U+,#�6�w��$�ٱ���֗W�eXw�.��O��P�/I�=�}q�<�V���5�c�I����7P9o!��f�|A���rқ �ފ&���.�5���^�\!��k��h��YuW}���S�d��:4��铇�!�lQ8��Y[�dzG�� �	-��MOHx��~Ѯֹ�UST]�J�LW�9R�n�a����������ӫ����5;9�Z}~(�"9�[�sm�ـ��L�|��@r/|�j~�XG[�V��hk��4�f�@G�&"y��֚��r� كY�Zǣ2 6tuz�{�VS)(�����λ@�;*���XB�v����͌K4�csV��~��ԥ��Y#X��������a�o��������a�f6��D�4½��6�/�JR����� ���@�]�0'����0d�q<�){W�~�7���R�f���c����� �:%Qw(�b������'�p��启+͌�
ur�c�^�������]�����x8����B �ASR����X����=/:ĺ':� �����/�q��#��)<� �	s,�5����d���X�\o�z�X����(�91���+���E�_��-��G�Թ�W��l0f����r�9�l�{�>��R��m�/y�m�q	�`	�9��y�v%��a��O�Y�����&�����'i	�D�y�nV�D�������� �T��Q�!/E]dԔ�mP'7�> ��J@�P��T���������+�[���K��������x��02��X���m���ѵ��ֿ�o�{����2��h�F�1��aC���� h�Ia��1&�͞�B#��� �Z�FA��
�1��E8�}5Q'�!yV@R#��;��mr� v^��2H��n�??�)^��?����b������aY�s֙8Zb3�E��J���f�ۀ��;���~f`�l	�jt�C��oN��FK��:W�KF�|�����~�rot���	fA��]&�N�6�?/n���K��D�-��Dpn]��tʿ�.|�:`,	(��Ģ�#^��Ws������B3�Yx�K{�2Qi�g$x��Y��C=�E�g��p"�e�P�<�%Oe'����]�Z�#B�n&@*��E���#T�N�����p�M&��^g���٢̹�va���k��� Xj�~���[iqm�V��3�N'�B6�m�3iK��x����FC�b&�y��u���D� ��%��l~���$���6?������_r.��9z��?�VZW(�H��c�apCS�N��{8�ܴ�����C���:ꏼ@�!V?PG R�xRf��E�_�׺��՗G��r"w�<�T. ����Ew����[�n�=�\W��1�����{�Q�����;��̽�-��)J�ٜi����.�V����v|#m����.��k�t�5�Q��S�έ����>x�Q��c���	�-\k��l��J?�����PǓ W�h���g*��O��|�RS	��≎���ա	c�<n�F\NmǸ��a�)8���#j�e���KT����φ��3��a������$=� �K��U�����"����)	����~Hs�K�j� a��h 
��w_o��O�c����븢�R�ߌ!sE���ۆ���o%[�ɉ~���3Fe*��{�@
�5.Ե�+hE�}��y���&�
:�f+�p+��ݢ����$\���1&F��C����*)�V�բؙ-�	��WE��r�I���������:�##w����?i���b���<���}��-��("�,�^x v"D�������9ظl���sD��oR}ـ%��UyJfL���W:�<��K!ZV�{�ɿ�������v�x/}su>��y%��''+Q�V��+D��Vʅ�\C� ���2;w:�j7��O�Ybp�m�C�,�ï��$�n�鋒�+�Q2�V������N�{�19�~q�)��7�U]Ů�M�~�:����(��13]���'n ?�B�)�H	��׳�_��Q��uEC�p�bR-F��-�� �0�R��+j�AJ1��>B�l���B%4���D�B7y#8�@օME�w�ӄ��d|�;��м'�:�W;���D�d��'uE�HO�4\i��V��J���_QۯL.���ީՕ�"g�����5<R*Ҟ�y[IHu�<ofU��6>t[��մ��P��$��U)�)�����:)�9��Ҿ
>:W꜊ARl�K.G�]��g�h��D�7z�m�w̋��gne�Rf���Ҕ|u�;�G�e���e���^9jӮ����:|��w��Z�J�.;��>�vp�^�	9��Rd�7��z��nJ�Yw+gƉm�l~fQ�"b�$�B{*a���e�R�\Ndc6�9��5$F)���T���1�_[K������>�:?��-����_�Oפ���"�he�#|����>p��*���業S��<���,j�"�g�]{�H46|�O�R|5K�Ӱ�5�����&v"�njj��?�{��Pܾ-��������{�}�Ch�h�)��2�&_ �x��p�^}m�y���VKx�V3
����w<�J���h�Wu.߀��R��ܓ���Պy��+�E��U|!1�+�H��lt�������ZծdcY�w-�?�J���rjzR諏��|?w�R�z�+,Ќd,�)!t��{$.l�B+,� �`������&TD��x�+N�'��?����I����IB�߽��f0����CH|<��G�����P����u^qz�:�W^�Ԍ3k:��\pO����0�v c���S��±va�����%�G{���9G��2s�N��n��T&�E6r��-'�i�ܑ�bN&0<,\ �g��1�+/��@��`P�� ?XR~\��ͫХ����vR�J2��i&F��9i�]�����L��G
8pz���g �����3kg�(�6��&c�*��(�WʾV��]wm��YEe�p���q\iB`�������AD{xz�z�@�t.�`x� /���0��`��	3�T�~S�1�F��>yt�����^IJ��m�Jqr~"��Be��Pq���x9�6�>2C�W7�� ӏ�Mm�A��/s�WK�v��=*�r�`��y!^HA]8W�vnԲg�%�n��7�9�o��bY����/�JF�Z�}xLB����׸�Z)xcW�<k[��g�����j�r�bh(ڍ��AZ�,��;x�!���7>��汶4�C��	q�Z���a�;i����q�D�u��r&R���zՀ�� 3��9�e����<��H�Ά:�D�	��
ٶ���x4�u~�?�>�H����[ �L�I\߄h�<p�P>�h��Q��2��;H�grfq� �C'�G��B�
7.R�}�ͤZUml�6���D���K�#e/������Q�G :"�|J��p���j��d�-TG�w���SP-�V\��Ö
NV���M�X�4	��
Ƈ�PfUi��q밽�$n�c���j���0`�]�?���d,p�o �{,Q�-��^��+%��8�(����ٿ�{ϰ��<�zH�%K�z�1�Ɠ$�p�q�*�ɩ�?C؁&�moMd�s�J�,}~߂�p䥐ln�~�2@{��՞��"o��Õ%�4�>Kqp�,+�8\L�h�V ߯���I��Ţd��[@��8�C�>���V�w�K����Ű��r�f���;r]� C�t�rOQ|'x�%کBٽ�(>����+˹
Lk�L�%`HvuwڬZ�l�mTZW@|��t�:�o�Ò?p��ji�|��o�__���4�r_7�����	lwqi���؝C۹��!�bc[-�(�?���k���p���+��>��+è����C�����Ä����P	�=w�B�=��a�g×<G�a&���~�]	������Q4���9#�lT}�r*J��o�|('G��n��<_�A;	w{.��cl,��w���,�¶]��ӫ�8��"�Mq)�P,����,����/�zg�������6��P?�N쯺v[�V�/g蠧ߋծ�dWz�ϼ��MF�����J���H�,���9V�r�C����0��>m��]�yC��D�0�P������>g%vLq�{O\��[�x�z��Op����������:)��ȅ�z=II�϶�nj�@���o�qZ��W�O�� d�4����^[��U����*n
^�i3�G~��(�G����lFb/�K�+�����;��0.u�2,���i��[b�&��㛘+t׆�4H�N�	`4q�=+S��"YeȦ��n� �>|�#�T'��r�E�X�ǁ��y��#ċPŲ2b�]@����#��<Z�t��x�b���S�����H�C��%m ���1~�"�b��S#��W\B����1"�ݷg�P�g@r��\0	a�W��f'�#IjLP���A9
yl��|Fk�� )q���[��#ә��O�P��j�cq�N�D�3�G�(�CjR7u�[2V���o�K\��е�ȗ��t��T<	��,�ǑAsY�?8y��������ɫ�� �`�\eT���#��%sA�5Gнh*`O���^Q��Lh�s�h��1l��M�: �j��^�)���)�Y�B� �p�H�A��g�#Y�]Ѧ78�0}i�|OhA_w/5i�)朒���(^�3����+���.��&�ۗ��Yo�jv/fH�\��b�Wt��
����2�e���n����^�n�ޤT��P�#�j}�,�Z��S���\�ɳe�R]�ȇU��^���$T�Xx��>
�U���=�����v�ž7܆>�V�y��Z��X]S�����~�)y�1a��"����������^
o�X���/�&蝍�J�w�Eϴ���1ߍ	��}4
bL� �*�H�X`�����sx bC�Y���x��*h���)��s���yw6�h8�aDͤue����g[lj���z)ES���q��W�.��Ġ�2L��$=_8D�s0&�c��l�X�U|�5p|/�_R Y��sDt�H�yÃ��'�r̥�UP���V�s��H�ٖ	{�s��-˘��z�t���]�%����'�`b�{��we�fl��2S�WU���38�-ª�a�agD�����@�T?�qPz����[m
B�;G��C_�.c��k�Fп#�Jv�,�m�j����Z2? H�"�J���z� �!@��������φ������S�2��iv�ؐ��P��7�%b9vP8��M`
n��@����L4�SG��Hds,��d��G+��'�ْ��z���kc���������V��{�G�݃r_?�nZ��&�V�M��띲�����Tn�=j�r��['����$��,?=�c�� �v�P�@�I�&.�~9�������8o�Q��)f(=q@]�U#��	j���p�|�C���۵���4��.&��n�ˡDVE�0I�x���(��*{�f�}�Z��u�"��f������nV���Ěg��ŨFm�ZJ��֓|EՊ'�9��Sk�.*O�z˿����[-�k������%"2��]ÅBl��=�q��PZ��j�<�㖁.�W�=��l���?ׁ���
qN��׉�ƀ���m]@����c�t�V�9�K��@=��1��knB���K�0[n|�Mxx��YH��Z�LQxY��:����}�&�.늈N]?��A�#v��}}&d�q����2N?G��^��M��[N
ui�p��x�4 �F��8����1����X�qP �����Zw�IEW�(tQt�-+M�Z�xO[i\�K3�'.+j��P3�//�]��0���]<�&�\!��%�0�ȳ��#���`�ft8�6�'*��ZT�=d�N�τF"Zk��^)�����ZK�!���N�?Э��x7��MX���'�G��ySي^O$�۔��|{H�b�4V��@���1>�Mu��|:��w��W�Y
��7�>��J��[���M���ە:�yt���!7\4T�G'�:(�ja��U6����^����ߍ��U:���wx3]��1�)߹?<�R=>�pټ�j�,!Y4��$ �
����E�=%�t!ѷ��WEk·��Q��L��6�cg�-u2��y��7�t��I�]�cDV,�S�1Bضa�pԓ�������dj���g����y�ψ~g� ���9�;v��-��z*�P�!�����x��R�X[��T�"W1�jt�\���<V��*��Pm�h��ϑR�;�����K���{���v�����D�t+��[i^��[���K������#�4z��CY��x�h u��q�$�\֠�<R�~ؕ`
��	f&��k�J���%���g���b{D��$�NY��وP$0^3��K��O��B��&��8bȭͿ��<?*����o�ʪ����D�E!K!,&�O���R\�?/�hwzS�'�����a�@����X�'~J�0S# ��t'e]�q"��$�Y�a-!Lj��W�S�Q0���X�Vv��<�P
rY�[4p)�#��v�-)���i��af��^�	�z�T4;X8)�.��K��<�|�~]�JZ����W瘶��7W��Ư��$a0�;#4���J��H���z�5�-����$f%�O��*ee[�W��s˗
��d����h)�n��=`;;���Nfq�{����`���X�{^�4�������f��}	(��FO`�
�߇q5|7�X�/��v�Tk�CBZ�W,�4eg�����jM�y�"Ne���	�t�J���z��CA�T�S{r7��P,hF>3�犡��p��3�pt�䈐���]֪5��N`�C*�-S�w�2���F�0���&s�Sά��s.����#���r�;��h&� ��]��vg�
�D�������2F�Nt9Щ2ԁK8'��u����K�w����v�~�J���mh�!�V�ɑ��Ԙ@5�j��K���V�"���r��05�^����3�*�\��RnVo�\	��W`%g\���C~{j���S��� s���g�q5�q�r^2��c��+�}��b�g��#5�N��(7_�������m��
�>��q�hl-�jPAA^��U���MmD�rBo0�sn'2����W�X>�s�~|!*�����A�^�Wċ'L��xI��,TB�"�׬�΃Ԛ�'������tD�*p��T�޹}WËǸ�I̔�	e��u7�gI��)M���8����������ۣ�/bL��>�H�W АF�Bl�2�?�V���f%/���_[22�&(��$~�k�޿ܧN�Y�.��fNmT�.4m���_�hy,���,�֜\�q{�FṬ����U����|1���$�yR�<�h��4�xb;ǂa�<^�~Ô&6$#����D�5%��p��DR��Ӆ�I���Y�͓�FA��@Z�o����>� �6�8^�ͤ���=���m!v���Pg�uI��M�,��9(��i)�	��b�Qq�0�)�YO���ωu����%��66���E���{�u9aȪ~�s������,b�n��mbV�8��HM�<�*�]��7�B(3�s��B��`�:�ñ��40E��j�s��������▃�B�4�	\w��4��n�5������;7�(�'=���rY��G���Yh��N�;qnݟ߿""s�f�v� L�H�^@��;6��<~�-X�K�5Qn
�nr�=�^�<q���	��aXr?��y������W���Cq��IAP:o'�4�y��l
I[����\>�/�Za�x3R�s]cR<k�����M���\i�c��G�Ni�R�N�Ӽ���y��{������u!�SX]�H�=[K�o���Ssv�o"p�,�cC���F�E�����S����ecU�`�����k:̧/��Zh7M����Pb�Cd�w�r��.�D�Ҧ�6ʾ(V6��m���(��wJ��d$nB-���k۔]��3��c�g�}�4��t�s�D�:7 ���\ �G�q�Ր1��n+���h�c��h��I�(�����>����G��<��s���S���&f�������	�W�$m��p�Q޵��?��]��q�>��l���C]�u�}U�s�WJ�k���i�����Q�੬׫�<Vj�v�C��;�d�9N�'�;��p��z��Qj�f�nY���%��̕��3������!Дa@��~�����qP�@�~ҺiQ;�z�lS DЇ���kSz���F� ��m~�(E|d��5�����5��q+\�rE�^ �D�U��)Y`IGJJz3�%�q�|`m�J�i�����M�3�G��G���t�4Aa毖�n���lm]n�	�()�<�,�.����DPI�Fã��I(e��U"�+�^:�ް�nVȗȣ�>l W*��G�F��$蓾h
Y[��S(�K!����ȥ�)a��� o�l��I�L����tX$iE��$��2��鵩WvTlCsJ-4k��_��Qu+��?T�?U���]�W��ǀ X���g�< �Oմɚ��A����������/A�yJ��H�nL>L��zg�ܻ�ڈ�^�$�]�M�X$s��uU��Xj��'���;�\���a������t�MVv+I1�xӯ���W6qvgS
�
�D�D�!}�Ќ�A��k�\���m��t��I��g�T�	'e궁���Po�}(��M�
mF�~��_�������'�rHfTT����k�S�+���fo��5�%�����?��
������u��%!���0�ڴ3����[=a*��S��Lv�O��\����^@�d¸���[��׏\��$��Ѣ��S��*l|���Y�<�1Q�fC��4�%&T@R�	����خ���b:j��}e �����������,ƥb�:ƬJI�Ua{@��]��7=�@��z��"�f�'��JA���0M߸�+q��Ҳ�~�]c6���x�Wb(v��fa���UF�)I��K<�d�v����
%}�{uk�\5���R��su\k?�N�N�j����)��Za;H������}�����TK�P�� @��%�4�/��e���(�$�I��������;yW\BZ��q^JjM/�W�"�����5"S�����D�'Z��G�$���$1F��5:Pۇ����	;,frE�B���kd)��~i�O�z4gˢ�a5�.��8��{���3����1x�]s�W"u&��k�%y>��2\��F����7���-�Ⱥ�E6��cw�♦�K`���H�-g!�P�$���FF�W�#��^��>��Ʃ&ތx巌����&!���9�M }���l��G�I�I@Z�<ǅ��Cb�n8Λg:~�H���:�m9�k:x���]=�1�Ô79�C�`2��_�c�������)��T��/Q�qX|5�=@y�b�E�����_*�م�a9��fB�4�Y'�As��QM��v9(�T�Y�g,-�zYG��Џo�Q�Jm]�I��"B�B{ ��b).>�ug`�i�X�S��} ��k��k�C�[��6�AnQ�j�=p���}�9[=s�d왮�,�Y7�mې��� �U����աI6��I�R�e�V�䣳�T�c�B��%�%�0�]_a�"�t�\���������ܨ��]�I?��4��+L񹺹�YD�oz���5Vc̕�����p���k�����lE�·7jO!���P�V��p��8~�ۡ6I�6���rJt�S�9��7��t�fC��I?!�����Y�s���÷xMB��o21�ܚ��]V��{�a(�a@A	)I�ba��9&f��T��
��.+�P�W��bG`�`�_^����YΘ��3��+{����jʜ��<�O-���~eJk�z��n���8�M�C<)�/��WѰ���=_s�Xzwے��xJ�@f5�jod`nŃK�d����'X� e�\��Y�!T����Y���.+��D�i�5�s?�j�22ӿy�myL4�I^_>^P�[�eyRdWƃ���F���9�	�4{t��D_�u+Ϗ���h��TrX�x�4®���:u��Ԛ|���׷�a=���ޕ`��/���]���"��J
�6��x�r" ����sZ�Y:��j�Q���,��VWV�HAY����#yp)[���4%�˯��J.i�)�9Ig!�̆�v��%�s	ݯ ��b�T�=#��_�V~���J�0�� ���!^��dI�ni���gU�zª+"M_�&���D:��]���1C��k������B"����p�� ��EY����&ߜ5���~<g���{oY"��/A�5�k��Jϙ���"	xb�4���!�zU�	��a���e��*��m��|4���h��"C$^�no|SqPJ�-�{ïp���CT!3�0��%a
�����Yqjy��Td�5���ª��y����z�7MyM��G,�Ӟ͟��35�2uH�X��#)#�D>2��{۹"��:��b�|�ҿ��W��>���� T�Kf3j>Aa�N�Gq%�2t0l�`h��|��_+�|����Z���zKN������/�P���z�2���Q�ѻj6k>�Ia����W�?���I�'��qB�c�s�Ֆ�y)@Ѻ�l��M���%q�@��3�Y�Ǘpe���`biC�g?�^@B�O�JS(�!B��<⋲F@f����Lu����2s�+ҭ�'��:U��Kd���2����>��$$�>;P�Z7Β�������np�oa��Y�]�؇̕R�4Bsh��զ����YK��J.�E�!��|s&���ҩK���kT}�wb9{���� *��8�8*z�IJ��WGQw� ���2{դ�S(+�ص�j���}+)0�DK�ʣI�M@��NK���OW���»���́\0��V݉�� XD	�_���dA('3N��?�c�	�pY�#㡶� �Fhd4��Me$Z76>��N��-��5{�mL} P�Q�cg5�����K{�s	W\��0U�K�8��
�"���P^�t���)Ǯ�pN�!S��y/V(�x>���C�`�l7�'QZ{�k4Z9�aƀZ-�
7�'���{�;��wަYG�)�IeNrq�G���x6;k'�`�' ���5rK6������BC�M::��KqGck������>4V�!�����?PlW����ti��V�[+���p������$���nU�y�R�{��'cA�]�j�x1@`*9�B�����";2���Ȣ�l.���+Ǯg�V��9�*��I�$��>?�����v�R��I�i�>5۹T����|b��n:����k��A�k�O�7�P��gم��B_�8X�[ƪk܏PXB�h�e�lR2`��Ղ�@�"��U?�	����L�%2-&�DgOݟv��{ )E%j��>d� u��x���XKl�M��ïehG�(����P�ON6���J��d�@��'h��)ݢ\���LD;���=z�3�M�)Ijb��H��x�]H��4��$���G0f���K`�5BFw]�W��1Y��\���cK�0w1�^�[���81���VW	�w\Q�ALI)P10{9��y����h
6%a� S	{�Y����urI��2�/�祟�&�.�Ij�&&�<�$I��'L\�_��'��s�=65�^c��ٲ�N��Vy��j�
�2K�ͤ���H�2SM$�!�PW�"c͔xw�߅G��'�A��6,u��.�!|P��Z#ò�Y�Y���Z>1`�s���$1C����?b�|��_$B��RTe��QηB�1�:2$�Q{G�ֽNw����ߝ��k҅�[�)��gL=E�>-�:z��zPԢY�>��>�����<?jg����l4��?x͡4�*+�Sr�[T�k9��������A��(	��Y���< E �p��F�q�� �U�zC��ԩl��s�/��FP��v8�9Hp���������ˮ�g޼�M����a/m��+\�?9�q�U�,�3̮1��a�	��u%a�����\�)I9�Hd#m�|�]�|�Sbg3�)�|ȝ�I���MX��)�����?��h�5e��)]z���D�R�Y�5�7I�;6����p��c�St�h]����~�ƅ��?H$�J6[ �<�aX����2����n|O����W��I�_˾��y��C�n�XV�1b�[G0�pw���ɀ�q;����&�#Jc-ii�ί�m?���AI
���w��䉌��-�-k��1ىX�
�w�T�FK;��(��b��3��G
���mM��OL~�G"۟���ͭm�,�D��4x��.R^�,`���.����nJ1һ7����8v��4&e;-L��k�\��"����d���nm	M�
:�كS�J*��M�����wMK{C�{p��AtB�C���Z{pIHIxb}�44�����؟*n��4�ԂFu|��w���R��U�{�xѓ��7�Y�O�.((W�l�N'M2@4���	���m(��9
�^��0c*
g0��ґL�|ʜ=��>�cj@��糭�.0*�I-��orAI|>�����Q2㹍�u+Z�Y.D;���w5�4c��ڴ})Ǽ![`�տ6,���At<v��XD�*N��2��d��7�ٝ��*��Iz�"d�� "���:�y��,�Yd+Jr}�G���`{�p�T�i �}��n`����Tót\//�xMf�u�3�v��G/�>�slH��d������Ь�7l��v��"��Y�/��x`�*�_�$A�듨g쐣��@d�j�c����k�������?R;�k�M�˂#������ �<=��M][��O��g�Jq�(+8��<��3Y���Tϩ[��'w�	[#���	Z[��D���`�0��rD[(�@���$��$b��ko��gpĨ� �N����}|��G�>�����N��J�(|���]�3�˨�p��:1�W�-j�}���ty�PyT>|�V������V2ϟ�FF_�$�h������y�b��y�L!�vƞ�T�T})NX����N��b�#����q-��Js Ys�)��:fy��8q�`��\s�6�L=�:���@`�w��D���������1]����������Ѻ0o�̳��6ۥN-z�h7�'��E?�?_X9ǨG�Ϙ�)_�D'|��E�I�_߇zB��a��W0�xYu���έ��P���/Q�T:��A_8J�F��w)	�Ze�d_�@&!���\6�1��GY�22cl�Ipgր�4�}Ѽ�=`c��wj8j��N��[�|��ߋ��+����:��H�(H��W�����4��ϻ�hZP���	�;��y$a������6(��"A�6#�u� *��ܤ�zz�\_p��U�b��N�!�,�0��½Pv��t�Uy�=J�)_��>׶j \�]X�t9/�йr��@(��";�'�Q	�)��5Z)���7)��l�Of['�V��X����GzzԴ���B��~�eV�-�˖U0*�&L���"�)����-�D&��明9������jAx��?l�\`�5{w?zۯj�,�#t��Ұ������l�ZA���������A�F��i��n-��X5冈��_E@"f�v,���+h�%䌎m�b0ޟe|f�����h�l�V
�BBd�bʪ���M߁��ܶE�j�&�Z�5�wBY=�;��	;������/�'��r`F�8|���df����`DT�Ȓ�?:�{b����Z����$��i�`���o��Q�i��cH�ӽ�c�&��R5.����o[��x�2�^�i#GT����NIC���>S;� �$���Y[���\Ij{���'J&��~<��8����8�яu�䇻����S��G��r�;M�A���P����	T�۹���7��K9�ż�uh-}WG��1Nc%�I˶2�>g5�ĚvD�>�C@Sy�f��'Go�3���b}b���5S�7(� p(�m�;�����H�1�Y^�Ptؓ�CG����W�LDt�o$=���P}�2��^y}n�ﮫG��q��V:5�=�:nO�y��9 �N���'u�N�ʃ��gQ�J�v��8(Mh�]��l����HT>-q����sKg5f���"��(0�x5p��4S!��x�'�-��T�i�S-8<,�GwmL�>?��@d��O�Us�_�n���·&�D�٩]O�,�h�#w-W`���2[^N"�j��y}��>R�X������T�s�ȸ=J��Q�}��;	!Դ(�G�`;��E����I0��Ƹ��El�[�@���Şv�����B�?��s�;/A��g���<T��ҁ�^����(�Ι!'�:��r+��v�c�g��e��߷�]Uڣ�n2n牄Z�Y�r�ӅWH�՚Н�Olp���1*��'y�BhױB�_�m��� ���-ߓ<4�eԵ���:~�F�nDK%WipN��r�	N������I[���/�'�A$�s�;�u�3[?i��gu�)oQ��}�z�ۧ�>"݈t?�D�WF���OK;��X�G)�B|6OE�_� T{�h�J��8I��:�9��U��_k}��#l�qVMtEt908�Y�9-�_LS�Ş :���h�]�u��x���dL~{��;͊����[����ʆ���W�1���rm&���X�T'zB�&:�RS��/FT�z%���K�,.��nG���Z2�<�>N2^���sB�RZY�Nd�c·�-F�sWxI�)��S��<v���%��{+ ��F�/���<�G(c�1��;��؛�*n
���<���c^\�ʰ�7��F��c��'O8	/�r��o9�z��D�D���#<�?���C�=70�g;�`�,0��N��[�r�]w�{�!ں\����駷]��k$�S�-���{S�0�����N��C�v���j�TP��-�mD>C�Z��tj*�X�*��D6����4a���ܧ�4�[G�դdE����Sǥ0��X�l>=��S`2n
�'���zU)�l$=�nms?�a�>��HK#P9Y�}�!1 �꧎��2fS�.rP��~n=�����U����wGdeL쓻�7�7�<��e ��0{Ka�@���oN�/��-��3��z|v�8X�a��(��0@1��6b�/B�K 5�ktK�o]��U��E&<�=xѱ��b��{�pO�bx@���e�{�������hH���	���V�HԖ�l�
�抨��&��F|����m̈́*Ip��"���őӚ���74�"�8��D���j��ʺ��e��_����ֈ �}�Sn9���Z��y+s%Zaa���1��sy��O��2����?���v�,RX�僂5<�)��q���T�\+$C���,F<2¶i��8�����_�܊5���J���{�o-���0/&�����yx��񄔩��r����R�b!����(�U�߁�~p�Ct���>e�jbK"d#�Vx�c%��X����,W�O�����|��4�H��)dA1i�`P�L�&���
�K��Τ���Q�%�/`�Qx�~���,2F�� �[W��&ћ����e�)�N2%)s��;b\�J@g֋��h���\1w�j�3I����[�-W�΃������4�!�B�^�n�g�,��_�p��O32f!q��{z�x�
�k�X���f/ �`����_~�H��SM�!�%�Dtb�,Om�N��^`�W����5P�����@���N1�`�r�@��Wiq���R�@e*���#i�,����t]$�����4�2Du�4 7�Jgo�3��hΔn8����{{�bL����#)mѧc�iY��������ԑ�>�'D�D��_5�w�X>'~n�T��q�<������~�J�q����L�����i2�ECx�� ��ְcC���z;1Q�V���̊���!m��gN�S��)�C왶x��_�i��6�L��X��L��:E�[��0/ر��YHW��xyɺ�7�d��dWh(����b�"Q8<j���EO�O�3u0�P2��B��Z��sCFi�w]Q�)ۋ	A�;ޑ�&Y��\�a�-�$\���q�m�_���>�U1>��kf��# ��5*L�/���bD������:<b��Y�k��p���%uV���@rȀ����ٷ��R�6��D�K|YأD�H�Z�pPǮ����L�*(�
���1����P� Zq�75��ԋ�?�F@Q
,I�=D�,�e��(�d|�IJ�/3�/�W\_��"��CZ�I9�PDLs�"eA����n��� 2�u�5��$�IU���E��/b� �c�j�:��kW�����V���)�?傋p#}�r��@r�O����RfZUe���)Y�T�2!�:�'�-�DYLԞa�uN,A���V�>�<�/�����nΝ�M9>�ɗ�<HmS'#�݀��̂�|2'^��g�?ä�ML���W�m��N ���t��ɶA&�����0��� |I�_�9���0�g�
Bզ��b��^��S�����bȶ!b��+6�c-�h���Ɲ,H�]ŗ��'�i�M�c	��(_|��	<�n�M�[�~�kW���n�c���U*b�)g)!W��!���R&��ě�?|@��g��^���#���찯���3JЩ5JW�����(���Qm}{y�u/8`^HU-��n�X�d{�a\�%�V�����8�pP�9_�^����a�H\$�%�3��S:�l��z���)X�����t�D�qLp�2\��&�����Z5v�sˢH�@����R�wҽ�Y�2_�-�6u}i���t�1Ӻ��c`AQ�v�r ��ѥBT�]-`aO�E�ٴ�Q�=��9����,��P�����}���z}Y�c
e�4�����3��=in�Vf��ڰ{c�~���z^�كC�g�_�#��1¾uc��?Σމ%y돥R���IH����\�����=�5T�[�i�R�&��
�'˥D�= xy��C��R+;�*f��O�+p!d�/8);�O��S��S�d�k�.>�Z�����fl�\�b��A��5)��G1��UFj�q�{�$e�LMR�ۤ;��Ksc��Q�_.u��E�S
�n�E�����?J8�/�5��u���颶��nĚC���g&�Q�1. �)�T{T�,�XIf|���ad������ל~¹NlV���;]wjd�D�" G�i��^�s�W�ʸF��"y~�Y�\���C��4NOZ#�<i���qg�:��v���Љ$�qQǀUA��-H��7��ӅZ��r��8�U���H[0������_B�8��V?�iU���M6��"]�^�A#Od��(w$�L�:;"����v�dA����^ǡS���4Y+�x-�['�O0q�7S�4��U�G�S�L9t�* آ�Ix��[,8���Г[(��a��u�~or�gS�.E��\,�C:v��C����|�*P01�ck�KI4�y���6F@�&�ΡՔ�ݵ~A+�nj!�`�����?6�ܧ��<�{07�����_+*#�j��Z$aEe�r�R�|�
�
�CM���0iFU�9]��rѡ�����tᒇ��Z}>6J{T(�'�֭��~����֛�u=�����n-���=�gsB��P��T���U�+ύK�(�\�h�%��3O�
;@������]p���c�fՃ��n�\h<K�+6��3il�0�`�8�(�����'����S��w f!�cK�gT6���f`l�?>�y���8/�6C���3p�
��P06���-�Y���C�+%+-!�b�u���a��T�B~�K�
5_O�_�oQu�#����c��6���p���t*3H�(��z�=�k���d�T�M���6E3�غ�[6�?O�rS'΋�/5�qY�J. > W�5�v
�
K��=�t�iB�֨��:�I+fD����C��
:n'!ަg�Yh��D�����ׁ�;/�B�@#��V������"c�&�M=||9���\�����S���A
ߒB��������B]��S�֯I�O�m �g�M@����ֵ�	M�.֌��o�Ȑ9�X�Å��:7��l4��^W�i�IV���?@@�ط3N�=��+[��;]�[�B�{q�0y�nqP�4�{�kh��|���F}Œ*!�:q#�>��5���Z����D~l:Cy���_����M<5�� `�|�:ޚ�t����7�H������_c0�l<&'v^<aA��RZUD�~�{I�A�OW8ay��?N�>t�S^=��"R͵��Ra������;�mg8��Q���Ͽ�%��D�Y�<d���b��JU���~ێ�	���]��?��1 �ȸ��oS�+ݨ�M�CV���!&���`�)����:^�\�o�x�{������| ��5)�6%馏X���NV����>�o>�����r���jgj�7��KQ����]˯V�|���l�k����Y���ա�Z���]��s6�C)��%f��Cn%��`�Q�A����r :v�Pu�t@{��T�����U
Sj-2���t�� ��mbw;�븃W��҆5�[����ޡ�V̫��<K���g`�|�}k�cy������d����@S[luFRܦ�6����U��NmӒ�]�S�?}U>�I��Ny��!S�x�RF,���oY��/��L!Ǥ8���I��ɒ�;�v��V����3M}�N��s��TP�=�T@-��v<0_������%��DTA+��h��]��>�Q�������L/���a��n{4|� �J ���+�/]Od��Ƿ�1��o)��Zt٬~9�k+��
V��l���!#�
����Q��pV�`$r��AX�)Ew�˂g�9�x����q����*��N v��Y<���/�T�ѥ�z,����"MD^�Gv�A�S�z)(9yҹ6[j Z���E��#�B���o?�ǀm)�<�����*.A�"���2YC#��cP�V���C$ڴ@�d�l5��0B�R�ԗ61v�i�f���#В�\%e5a����k��*��5��Y�Ќyh[��/(�p�xGǵueZ�-�xr�ۤ�3r�O߾!��'y�\��[~Y��@!,5���fJK�p��D�y�t	��ͻ����j�)[�Ǚ�߅�^����,�Y0G�2ˁ��?U6y��
���`��}$s��G�+�ي�Jo��m��ĽR�ar-=�g�}�������s�-�������( �s*�ӑY\�k筶x�e�J��{d�Cخ��}����E��6
���c	bl�r���`^X$\?�Z�X�ŉak)�8�%�sl�i�/�9���a��h�س���Y	���Lߑ ��U{��	���b��t�(���[N}��gq�+
vٮ��2��B�7m�svf���W��4��"��&�-	�n�&"���Ɔ�!���\�X�� 8�D�s�O$P`P�g݄�_:���j�t�@�e�	,�Ss�r4�P��d	_~��v�:��|B݈$7Dj�<��|8U��O�g��~�����@�T�Q�$G�_5��eu B�{��ڙz&l@M���b��Q�j�:������A���r�w�͉ܔ����G�2�f�����5��>�s+b� an�{��w�`�jY�6����QQz�[�����0i�����\��ȂT��w���D�K���2��z)i�6Iy_	���͆{��6� �ه_Iψv	L��qӮ�	�}�6s��� J�z��]��<����p��WmN���
e\	Y<�}�M��-�Kהo��hM�vݠN���M]�y��f�Ca���ϿNSXW���_wg�Γ��0���A8������u9a	Ȫ�����cQ�P�OY�d0�*�֊
:��As8�_$��*=���#H��^�0���	.B��� kw ��υ���'F:�"�GJU<vk�����$W6�h�{GR�UEi�'��ܢ5N�H��C;���V�5��)|`!��	�۴�<gT�F��S��L��遲������5wN�ӫ���c�_IfQ�Xݮ)� JI�l�]�i���dlR`��&�D��D_�,Fa;�o�oK�\�+�,�d�SJ�B�=����m�@:ܾ��QQ���]��܉�u]����HB��,쐪�B�uټ(�߻��3��d?ǚ)�cuφ2?`�s�ۜ�P䟈YoX/��ӏ�`�(i�a��:������D���G�^�B/��mh��2iAk�gĊ���}-���w��e�S�^
߃�|��*�93���jI���u�
]��A[+��Jw|�Y�nd��E��������td;��ӖJ}�ڈp��0C�ޔ�t�P���dN#o�X�*(�Us�Ԏ(�>a�-kG� >|�+9�;��:�da���|-��q��z�
���@V*��	#��F��6Ȁ�մ�Y4�f�x�2T �t��\:�U�7�ӣ=�D���s�O���%;�;�![�䄮�k�DA*���2�xi����`{T�0`����m��Z�ai3�/,T��W��Pk@�"�=ȯ�I>_=sIHC{ZK�F����n�K��i $lCj���2"�����S|2�eݾ��/�V�u����\Nv�{:I�Ds���Dd��y�����	����g<90a�A�ٚݦx�%'XQ�� _d����d�4�Ӆ�p?tʖ��P���|  f�CD`m�d��蒎V��s�������w�6��#x:e��h�9�Y�GyW�J�LiY��1-ꍹ����ј���<�m�\�IH�4���1��xU��g:�D��i��t��ص�D!6�귰�#�c�*d�z�i��
�53�Y��f�O �j�j¨R&HU��A6�
�	c����~�ϥ|p���à����D�������}�3Auc���"ﺔ��|#�7q�*�������* I�w��ls�� ��[��0��V�b��[~j��&:��r��BQ�i�����Wr
u�[G(��40s�VE�g4<KhJ@V�37>mIS� tz�{4���؂�{��Nl���=ӎ���e?����̨<�@Z�-:�e�/I�SQi�km�h}��w��ЄP�Iv�$ư��S��3�	�j�_�]�#r����?�4i�B�s�������-@Uc�kS��e�3�s����020��U�'�07����1�tE��H!ŏ��p =��'�7>�6���M�J �3�sƳ�)�i:x�c�ɍ������A�����8p��H8M���
%x�yB���Ln]�7�V0�È7�w�Lj��6V8���%�[N��2˜Z������$�b�[�Þ��up���\c(��.ޱ�K�'G,m|��Q���~)�B�Ge9&��/r��r����1�,��4�\�n
���C����\��]	����jl_��hqP��E���?o��s�a4�X�Jo&��}�T�V�AVe���xۼ	��P��o\?��(J��E��3�Q�߯�=9æ�G�b����>���X|S�A_�*8x	��p����W�����&��=��Q��rcs2G�������w ̉�w��,�zt�5oGeהŤ����Vt���X���r4�@?��#����Kg����zG'[��rp�/�ӎ��bԖ��+����3�,%}�K��*yγ���_�����&��}�`��(˭�a�=y��4Q]����[(�)G-��R����kc�y���� o �.�ՋK?G�9���g��1�Ή���� R[�z*X㐃�I,i���~R�
s��?�S�?��{z,�Ղ�N�a"d82[��x�|�"�Ҭt��e"(�91���@@�{F�Y�M!��,��
�]���`������uw|&JK����|���D�������([��#�;2f����tt��ǹ��'���F(�:�awك�ȿ��P$�&���0{D�K��u{vi �0�樂Zv�a����s�&(Ș-֠�3Jl^K�*��FJ� ��/��wʼ�=c0�������UX^��:2�-r.�����8��Ԕ���')J�C�HW����|����pA!!��Զ�z��B�GO�P���t�}I4yg1@�bdd% Gfi��!��P�nCG{������?%7/�xp^S�/»�j�`�?ĖS�`��~��uڤ��T�"� ��H��F-�f���,���3[o���}��}R���h�Y"��4I��;�~�8d�h�mٯ��$їP}�Me�<��-��%=M��4�t�_]�]Y:M�a���-�K��[��9������k��#B��(���_�\��������G&�
࡟g�1��,�F�l�,R��.��m8�lL�ʘ��.ɛ�9����+G��UBEK�ַ��4���/���7x=���o���sc��Y.�$���l�bP�℺�\�$[nI�`ZDƐ���J�M�
�,�bjB��G�3��+Ĕ��l� ��`]��x��b��0ᕕ�h�5��P���H{�}� �"�-Ժ��_$�ʒQ��N��N����(WI�:>�'%�l;SL#�I��R�u�[�;]V��+�e�>��~f�d<�vW����R�;��-w�n�u���Ě�Bp�:^�(�����3�H�2k�<���t9�2^.Q��./�FP�"��GW0=��i�E��ln����c��ѧ3e)J|��yu���L��K��YB�)�����ց�B
�$��% ��9)�@Am=6�@���z!c�*\� Ƒ]L>��
����X#j[rI�
�6�-
��p�C�6������m��J��r�|�s���?��Aw�̿�ډf�<v*~��e�z�F��{�3�%�+�X^�X�
f+��>�ce,SRh� \���wE��I�����M�&�]��v�4GS���n߳Χ,/�]P�E@��I�^�z2�;B��L+�=���a)3Y:YS����+��-�e���K�y��ر��I���`�8~M0��׈���I3	�Q�t�G��n�<��Y���e��8�,��Ʌ��=��_lH�ks)�ӽ�i�󈭭`��J�Ӓ��qz=1�߅V��v���s�5���ZdU8Z���<8��#�W&zP轋!���<D��?�MገM8��4�[,P����e�w�$��/=������<;15,+5QX!C�������E�'eg��Z�V��6P�ֵ�;��z'��]8�S�~?���*������΋yJ�r��z����$��*>�;�<���'�L	������1t ��1-K#7�Lt��[��X���U"��Յ�;��TH��,���j���O���RHox�� c���J���!I?S�_�SGEY��=��������x�J��o�)���w${_k,K9���dr7#�b�Gk�U��v�E�P�s����=��~Æ"�ڐ'��t�	���Zl�Y�"�l�\r�S��{Y]�B&F.��p���Ĳ�r�&}>�A�n�̢TE����w 6ɮ��p�˯.AT��>dfg7S��𝨦>��M��������M`1���~��݄�	�UYiW�ܥ �U���n�u�N?��|�e#���x�{p��*&��2�?pI��P&�մ��

�ݭ���|b=p�n\k��C���E��)�x�lqP����r���K�5�:I�?��8�3������~��~��a�}K{�	v�	3�nP,�0��])�F �M��{���!�D��š��5f����k�i(����Zזf²�r�lj�~�9�����q����(~��������ғB։X�ΜW#���>�_̃�9*q��N��S����y���s'"0�$f��H]� q� ���A����\	)B��a2�E�0*�j<�Y:�0����C.ɝd��d�Z�3?�������e(&��"�r���,��H�ĝu]w���W4�{�Xޚ���������jy;�p��� �XL�{:)bE�LN�b�d^��54��s�
c����e;�Qo@mA�G9)L�[gT�?�^��B�����s�i*FUD*����*$mD�%i�Ė�/�ލ$C[�rᓮ�)���W��Â��
p��0��*dj���f�G�}�pV+���%���ϟ�U��vg,y�Iw���=k�4�d*���Z��߅vE�A>3[b7`�;��KIX�߽	C�9|�$,X�ű�Lͨ���~�����Eͷ+���S'X���nc1��q�������D��3��\�>6V�B�J{���At��q�B�B��(��#N2ѰMA�`�h�Ux���^�d\�����c���E f��p�,E�	p�BSHO��Ynfϑ�0�5V�L�X~-G'�ֈMq��e�^��P�od��{Փ��!M�s�-��s5b�/fk��r@O��eB��.8"�nΦ|� "�q�d�0� �b��
V�Ba��Ŀ6)����M�?|����J�+�M���ֵm�B�YM���f��7�e� i��S�6�z�Ž��\x.��)��l��o�n;��B����hz6A�ar��+v\=O�V�IQI�/ ����!��GK�ΰi!����q-� �V�6d�{��Ȳ����5��ҭHc�~������Eϲ�ۉ��9t�z��%/�F`R4��*��1E�5�ŉ���e���AZ���ݏ�VVE:O
4��$	�Ak��7�ڧ�3�m#�h@�����@噲�XnAfa�Mw��L���%vt���҃P;�vp��"�n��e��+��X���z߿��֖�rv��U�v��$��S�JF	P�e�����H�~��k�
���B8;����*+_�XL�j$�B���f3d!((9+�Q�:}�O��3�P�$��
'Ƹ�b���o�/��B hP���du�0/��Ӻe,���=��01�4�-̋�@��t����Mi}#G�
ح[�La#�/�S�!9���]@�;>�,ɟ>��e}2?�Ǯ�E��b���0S}
u�j�&M.�p�%y�4�3��U=�+����Kk����!F;�^�|7����q
�C���q�_�8;�d�o��IύX�}���Є�!r�\��O<z��D���<}JJ���?'�H��d�e[�Ab��(��=���[U������9+^�v*�"L��S�;_W�A$l��v�w���Y^��>ӹ_ c���-��2���TSEb�f&��2z�(H,�ng3m[���|�=K��<Y1���&��hSN|���AkdA���/��!�*���OY.X����A��\�ڂ#��9q���c�5|�ƽ@�[�R�Ú]��D�������h�sݶ��k����K"cC����2�{�~)�Ho
���Ƿt9�a�A F��IS�e��	�O��>��4�w)ٵ��Rt����C�10=�wWg�f�#�"��{�tw�i��zR��az�*T.�{}|ń#�Tg}}�ב���Rt���R��^\�c�9sӺ�p*�GZy�)�q��^)���ю�&��`�a�,EG��M%�ϵ����'��y��h�SlP��-�y�� ����{?�b c*�P�� |5t�������C�D<y8 �����$\j�-��)L;.JZ.l� ��j�i,��$�]��}t���X�3U��qk�
_Zۢ��H��6�cE��8�a�<緅_U��Ur"b�Fը�L��-��6-�s�qXK�;�Hد���A�M��)}�˒�)��N����_�e�}�;$��T-ܟ�%C]�RnO�����}����T!Pا�a�ع�އ�4����+�>���2�H�T4��?pSG�Fإ�x�o+��~}�Ъ��NLt��^�������\%7�d� G9��6�������&�q�S_œ�c|��>}�~�]W�s���i,�ǥo��:e���eUUނ5WFn��Q-��5�X���0<�i <��t�#�46o��.�a�{I�'>t�'�6�je� ��� �v�?��qeҐ��WŭM����d�v�ԥ�JbP��zֵ���#�ɪ���Q��R0�?�Be?�`Sؾ��S6��w*@O�o��	r�R�;���y��ba/��-!���+Erǥ�w���Pw�LVF�h�_�T|������_�"�`�X���NPW��Y֝�&1�'{_��~}H��'�s��1Lm����Ʃ�iIH�O���J��D��g1�ܞn�/���VB�Gg�#t���>�r�sD�>�-q�j�XR�߷	s�6̯YJ�)Wj��.��Rr�)t��Ÿ��K�	"h����٥���?a��Nd'E��c��Y[��{�����)}�(���Z�>}^Ĺ��`��7/J����z�X\,�,E'��Y�2S�	��_��DL[f���
�`������h�&�Cu���|8"�31�R=�	�7�F@XИ�Z��e'f�`V����༫D����Je!S���~�m0�Tr��O�`�K̔���}4�����<QZ��~F~��'h���@�!������d;�Np͘�K0�&w@)dfEvh�W����bS:7%Z��0�����%��Q�F��l�g�ØH�D�a�Rs����hU��1X[	� �k_)7BnM�Xj���Tqq%n�>ޅ�[bT�$&�\6w~�v�Z$r�gP,�Ҙ��U7h%Sn���Nh���
�b�8���r��\��:��y�!�O�s���~���2��6�B��I����b>u�EΚ��G����������*�a��
LB������~kL�����]-��4��	�\�݆G�z� ��@]?��%]�Rx�����h��dT7�*3�}#�g+��-�oM���(�d���3$��J[��I���`m�Nv3�*�"u[R��"����ݡ�9��$o0��y����u��@��Ɇ/F.��d�\��1dJ#n��n�����-��ٺn����x�뿚�{�1���t�	�$$<{7�w���wr�ݩHB�͋�Ӓ?�8�z�`�N��<&nt>�[E	�a{b��@.VO�f��x���7 �6%�k���p����pݡ��?��Ya"���if�������.7;���i[mk�&\�B��Z��C\��u�d�¨K�������w�T�E5�
N=�������+�Sj&�U���pĢ�W����>)8?�?��T��yh�M zi��$�IL�$�����L��q�dj�˥�2ݴ�I[^:NkV#w�"`!ix�Ĵ�.����S��D҈�Ϸ�zEJ��b���?F]����#�?�oD����I�dV k�#;W7�$R>m�*_���uA�]PL	�H�rC'�y������D��ghҩzǥtyZ�-
��f~8�@��$YsV�?�u��x |x�����ñR$ ��9�0�0"E���Ǒcf`�b�M::�G0v��]�M �7�u8�޸O/b�ξ�e3:S-XCVi?w���#iBK�`�C_5�ȗ�~n坓���e���:�>��KJ�N�r�22g��W;��+��s��	�D��Zg=]"�2��k�S 3'�a�t�"��b�R��N����d麱y?}��]�I���ǰkIb=p�wۜ���+�_XJ=u����yd�?�.,���B��.Y2����Jă*�W��h>��c�kӥn� �3]�8���8(#׈s�;;K����oPU�$�U(x���P<j��/rR�?� ���q/n���(���-����\�W[D|U������V$@��V$l����T��ų�!(�]�NKx�����A��Aإ|e+���G��Q������������X�-]��l��Ѽ�x�/�������w���4�[��m��Ȑp��m�=�+_�GlsOEY�����|Yc��ښ��u+��%��g�T��6�hg��P�IX�p����H3V g��'�~?�i�����K��c�d7s7(��KG�Z"T�;ۼӗȰNM�����Y}����^�\���ĩ�+T%M�2W!O��f�8~ K��4� ��xV���aA���BrU��F/��LM۳�i�m�r�)�}��&�hS���[�r����YVZ.��6 ���Y�������q�^Pt�qRY���*Z ӛ��~&<���eܑr��`���lm���5Wr�o4@έ7�����?�i�E�+s�- �c6u���:�3|mcòR���"#�=��!��4)}�F���GX�utM� ��U�9c��h2TT2R�L���a��qV0T�SF	���w��'���*�L8>F��/�O6Mũ�]x��kN���Tl�B�UJ\o�f Y�&�����P(�9����s랃�����pΆ�@��i�7e�T�4�Cg���Cu��(f�`��n~+�����L��s�]�[���$a�����U�ם�l/�*�I��I�w���Tv6�Y�L`�V#eQ�]�� Iʨɥ6��/�@rp�M��tY�#��@�3Z�d@ؐ�v�r��&_#wFx�D���C�Sp¦�����N��X�k�����E쑰�3++a;�HT7Z��b��ʨ�S0��-U�����j�+��r��ƹ��{PG��#_�y�2��R&Sw���L� $�o��HG0����Q��1̵^�z�6&��Ҹ��;U�*p��oKd�.}��=�x���s�&Ѳ+w
@`ZE;����bVgp��
 �����CrQ�R�a&F5J�p�x����6�spV&��]#���d>�� p�`��0�sx��G�P�(:�Eg@�N.�g=m}�J������	T�v�g��l� ���I����7i@�%��&�oFYI=��C`��Ge ��St��1��0(�W��
� '�l�AJ&+pe,������\��ɫ�Cݓ`�_��<��y�Q̂�����M:ekZ��K�S�\��-.��R&r'����U��Ә7҇yE����`�`���@۷��>?^S�W4[���Y~�I ��1~�~�aK-�`����I�z;�v5�/�� ���f45�͠�{(ׂ�CF,�p��FO���-.;�Y MnS���r ��3b�K�n��.�[�#c4b����/��Sݛ�l�De/`_g�mtH���|R�t9Ś�L\�s䢹�Ӯ�P-�yO����~F�)�=9Y�L�	��oэ�^�T%�P!^�c|���}����\�a�r�e�b@�>�o+�	�a%�#e��ik�}X������WJ�j�w&���9'�Vi���c	���v��E,�3����� �X�.� �d�f���5u�E�]��Rj��x��fV,�x����J���~|6�9����B]p��Ĵ�JO����$����HM�r\����*�o���}�rr�cJ!��I��5����{�����5";}��-�Y�V Yub.�C��l��D��+�q��~x���G��)��#ȝ������s�\����<�h|�/@�"@��uD����}��`l�9���q�q�-3�u m�wW��"4�>.�#_���&}Ҫ��$��ֵ�g�i�9����u�B�ysV����VZ�6qx�]q��	��G�:�eg�����>���}-�=�h�8h�u�d�|e�XdB�.���p�6)4�h"^�ȶik��e�_�9��z��T��Zkׄ�Ք��x���r��X���p�S���ٵ�!ҿH�j��n/9��db5|4�e�4����L��/Q>@&��)7����n��xf��\RID/;b95=���3օO�U��2pHJ�
��AEg�;�*:�t*�L�Y�V<�k���q�|��>GX�f�L�악��$�x7��z�ڠ.��>��K2-h�z J�PDn� �F�.KFҊŧ(� \��~*�sY���˟?'|��Ŭ)]y��A����RL$� �H0�{�y[��w#fK[ �3c���$�G����(���3Bζ;E1����;��BY3���x����ӛ!�9~��4�D$ ���2�D��;���j<H�6��y���"ł"�`���λ����zbp��.^AG�C,{"G/I^�$�/���3�J.� ��]M�XV++$�������r��^��lu���J�P��j�fԖjF�߹����1��%���Sŏi��8���2��S`IB�ѾyWu�ަ3������,���5���V+"|�m���ͺ��mH�7g�s���j�Uv�\S�q��neP�tOd#=x�4�x.�M�8|���D{<��W�B�Q}���rt�aA�pE��Zj�����8��s�{T����\۰g�":�<%��>c�=�"����<M��!�PC���4_�\8�EW�a�u��Z\�˙�J��	=�o��E�rOy2)�6�ij�O�n��{q%�y���4:���S�]/�&���j"s`��^�7`�W��� �Ho?vZ8�=nlԜ$Z`�`�߇z/\����M�Z ړ~��( ���� BVWC�� ҫ#�����ۍ��������T�����B�3����H������ ���.�E��������>[K2��lb+��:��6��6�>���G��Q��Vg�X��ځ�ט��յ�P{�#0�����v���q]\0��Ҡ*���.8W��fW��@�P{9&(���,[`���Pj��ϝ���i2��sm�duk۷-�k��<��-A��Ĭӿ�B�+gȿ��"�D���n�h��@��m=Y*�LT�������w���.��`��$y�?��U��֮��ᬯ�\�W�z���.��<ɋ�ɼu�Y[EjKǜ�`���<$;Hmw��p� PJ�I��Ԏ�_���W	)D�������'?�����H�8V���k̛wP��^f�&?��*ϖ�*�9H6�o��G�;��7���tm?M|�xʚ v��s���hp�}��Qٝ�,ǅs��ߠ�	��>�'��/�Q@ͩ����* �a,���"��3ȹ]I���ybI�{����{X9�;��}�E�DS$�Ί�?����@@����Ŗ����j��(e�<`,"4Tj��',QU�r>u�T��/=�>ʛDQc�������z��v�ͻ���[D%{�Bv� �bA
M9��v�3�g�,Js�_a7�}c��v�^Ku���0���L��\�d��~R�M���yx�=Y��33���[ְi���뵘.���c�Z0���ѓl�љ-0l��َjh2͚=�f�liu�D�k�^:��Iz��u�v�"����ȧ `�iL�a���mrB<�TS�Xi��[�<� 5��� ����6��nҬKm��	`⩜�������W_һ}��Wm�ǛGGҦ�g$Î
�;~�UDHI�
m'��~3׬���%� s���u-�
i-�h�:�>�����R�pM
?��䂕��|�����9���</H�>�,&�O��n��.�\1����2k�"�e�PH�8�u���4mi4*p��a��f�_��c�I0�y㗈
�o���� 	]G,��������Gp�ts��wʷ=��\!'H�>���$���	�V�Y�|J1�x](�� ���K�W�1��q��вf0RMV����$�����p��Ϙ�umW�"|\E)�K�s��z.�%/|\���J����I���;�N�m���&��	_BV�ݜ렼�B��
}��t��W3�vdo�K��<�6r w^"2�#!9�ĕG˨.�q)r�o���>�=�Cl@�*1�,GlW܂��+4�?E�v@�Wf���j���g� G�S����½Ք���n��cLu/�e�Z����D�jl�W�!�ʕX�\k)Q��N
����;_���7B��p�B���s�6�U'C���r=*�<FF����۴'j����Љ����&�hn8)K��`��"��!4zl�y��;B=,���K�Da�Z���k\�Kj��f��]��AdO<6��(�i����<����DK`��,q��o�_̗ۿ��z��:��S+�6��\Y1��l�e����z�[�Q�ѫ�N?E�<e>>E �,��z;:�wr$���R�M�՝��QR��/����%�ųE�>�u{�-a>�k*C־�J�ʃ�L���v�@��&��J��Q69�ȥ�V��MZ�-y'��⇡��:�x�C9rU䉧��/��|m�Ǖ�����<�"
\=U��e�<���8���A ���`���7,m����^�Q�E�C҉��d9 =�d�O�c�)�b��;������*����Vf��&�ǣ�?b���Q��cc�m1{z���n��~���O�;��Ǥ@A�20X�a�4�ùY��s@��{��gOHez:%G��gd��j�m`�@$Z�d?]r�
���{z8գ�A���LL+���u�g�������D���m*�17��LX��>�s��zS`�]���|�FT�,}AR&9��2(��h(�O�>�Sȃ�������'�W��ǳ_��L�AT����,e.m���"8�����e�݃r��o�moRQ���vb͖w����^7�M c���TY���aq���j4��,���f8����eAe1��T��Eڳ�m�d,ȫfN\�}3W��%0���_Il�c�k��qkS@�,���mCR��(�n���js_��,ɸ���`���wOl�U��푘"��q0�Ւj�*���5ŏ�(��UG��M2u7員�ռ����^8M�hS�g�%���W¦��;CR�Sd<�,�����"�t�7rڙ!zk���Y��	U�⋯/>����T��\���d����DdSx���z�"�C�Er�0ޯ�ѿ��4�m�첉9��\�@�����W���`и�j#��B�ӤR	�T�"g���j��a�? �m���\Fd�BY�+u��V6g��ht<�%C���o}?}�n�J��b1m�����?��)�Rg=!�K,xW;���h�2I���u� $`H�&��ǲ�O�����y����4vm�3)_�0A���S���)�(�^ANI���ۤ8�+ �d'Xӫc$�K��B����fk��D��}c � /	�e5��2΀i��ّ�-9� D�nX6AJ�c������J����l��M��8xk;�fD�:ToVM�g��Σ��
�}�AlJE���i�J�z��[�����#
��K;I��Sq[�7	����[>!]�H��+�E��L���������e��F��z�A�sH�����Jz{��!g��Ps�v��j�����%�"����K�f"�W]�/���K��Omj�җ(�hO� (�[T�Z���h,M��������M �;�&0~�װ�_��Kã�G�I}{�v�dMv�<ŷҷ�W+��~ErRD�l�{}�2��4\֒��v>S���-H�j݉�C�[X$��n^�w��<�0����#a��9��Dn<��Q���9xx{Ns0+��$���	��� ����9)9��&�d���Di�Cv2h�|o@�`H���$�lR�w��i
���|ؓ�?��Tn5�_�k��7����+����yqm������-�LQ��y�[f�&h�9U�j��_�K~+{���h�'4��[�7�._������T�qn�F=VƗ*g��A�����{P�Q�mjn2�"�)6V�q �KN���FH���GM�-7�e�R�������Tdxa	�Xq�(&�w�y� d	n�vs��A�q�^�M�E{�o��� ����gk�X9i���ϊ�'E2�U�l��s��n��7�N��07���!v,�=Ǜj���b�$)Jq[6P���xҡ�H�\�Ts���d���@�#4''��	�6�Zo��k�C�IlY���h́�N$Fr���V��@�J��uY`4���.��ۢ���O�,�w	Ǫay��-�sQ'u���%Tb�Cѥ��:��,x�����j��R!;�)h),H�R�Y����SM�����39���r�@�|�5׵,���v}�.�A��	�p9�C�"?��k�t֧��ܽ<sj!�0؅p��0�s���2r]3�a�����X1@��lؐsrL>o�S��h�xH.�IB�;i x��F��4.�;���{�M2d��e5�^mP5܄.'��B۠Dc�>�6G�A�H�s�z�y����}��Mhk+tcU8'xWH��d:��i^����|�F�լ�+��8�$#�e������U�U�ZFE�`w.a���C杭�ɞJ�N;�5]Y��1�L��1��T��|ol�/')G�����?mS��ղ:n�M����̓�B�Ĺ�i�N���|��CV ��O��w��lU
�JL�΢;��>[�'!R����p�,�<y
�LR@����\t!�{��c)ȇ�l���b�.G���!����M0@�L�xd���$���QyH��걢��O;En��2}���#�$*�A%΂��c��R��?�O�Y/��}I}*��C�O���^�mwlhb�e��7��y�����'J@�^Kۑ֒ka���ݭ]��� E��$oq��4�x&�A��G<ɍn�I;��'�D���~/\���A���g<mt')Y���P���ow�-�$p����NHf?�������)^����������fQ�g�aT�Gi=!��)�-�5l�<����qK�Y�L,�3�T���
4s��[������QDg�<�h��4����ۑ� ��ܞ���F4^��d-9n4&<�����@6����1��+�b|�CK5��{7��ˏ��5�GF���]�1w2���� 1��xYC���c��9 �Y$m�,֯��Gd'	��4g{�1��@�A�+4�b��rP�Xc%�+ 鱔�� ���>���I�:������wXSUس���j�f��C��y�τ�ֽJ�tv���jC֢��5�j)�A�qZ��O�k�%��?�~@*v>{`��>��r�"F3-�Lܧ�$��겅Gf��Cl��df�V�'�3���ԳXj�ĚP�ꘝ��9M���4���4]Z� �rZ� �ƴ���e.��ΰ��PH�5ܖw���f�2������>��+���>ۉf^r:�'�7���T�e�{��\ɾQ�CHБ��O�'�j��mx>/�:�&VUp����.c����ԋ[L�SJT�2Z��Ꝝvϵ�֤xX3������Rt�Q8�z�]�����Ȓ�(�Lv����G������s�o�l�ȼtG�X�/�'*.�1��(���B��3x'(��^�@�Q�+��UB��G�Hi}�z$*�2���a�I�]^������ܨ��=?l����M���2+���	z�һ����x���<.�9�<��!�K�/�kdO����ɌL�0%3z#��~v�Q{�[�!��z�/���c���=�ã%[)����|!}�^2��� �ġ��y#CfȢ��Q�6B�x�E�˶��eU����K�kw>��_�h�|7��/��vA_��Wi�}n��GeM^A���¼L�A��w�b<>��;U�O/mn	�B���d�N�ş������@]AH��1�X�������� z\5��<�cI��,�4�ݢ�یd+��x�"�#<=9FJK�9$;-Ĥ� �j��{ψe�ל� �t� �GlT��OhD�U_�9�R�L^v�;c���jb&g;���͒�-&H��A8�aG�p�|+e^�������4�PN��قa*���O�ǘm~ �X �d�:�4��V��[�1��yܪ��S�%����_OA�Nd8��;�:�0����YD06W�l�gW���-"�U�-Re-�:+����o�Jg����̛he-���9|[�e>x�	�د�{Z����q.�k�)Y[�@�yD�����ҟ��~�*�����Q{r�0<15Tq��&K��z��l)P�٫��o�	�
-�O1G���N��ʉ�3ǅ�����ճ�\�K[*�	�Kd�qɅ��ە������R�=��2C!<�6���0�Z��fٞZ�彋WVКc��}ֺl�@��L��ܘϕ��x��%�k�AU���İj�48�KO���J�.39:i|���I��4�Wy�z8�BF����<�u�x"�=,	sYJ�Kl.m�L��dSX�(��z�&:�e^�?�S�R��w���c�}�,�"��9��@�=6�������3�w�4��G���t��������U�;S3zg���J|0g}�}��vK��r�e��xRۂ�e�s��U�6�i*6z4͚&����
��֤�:t��H$��3�O�����JB$O���� �2�e�,]�`�.��n9øs��d�isv��R�Ho�fm8A81ú4���1��B��ü�5���x��ԇ��@�L�h�O�8�锶���2â%	���(�`*����jGV���˾MI�]�`�X�8Ƶ1W��u��R���I8���j��v�~�̨��\�X���1=�p�O����ȹ�C�;~���X�=G���M�wM��/�7T!n'i���|�'�)\�h���#���R7B8��<_� �h0Р�"F�НP���b���vs�s�	�#.���K�D��uB��U{���0�y�������i`:%�L��>Nꆴ��t.���.,p�bp��<�K�Qit��#�����[��N�T;�_�Ìɼ��a�{�[n7-�氜�L
c\���y'���xٿb��`��t�����RDkBc�S�2��$����	���p�] ����c����OiR�vn�p	��O�1�<}�^5[��}Z/�5��?{.�#��ƒ�Z�E^��l&�ĭ��Q|
�H�am�$;0=MUN���`��ʋHbX^���r>�O�<�@�'g�@g-��8F�v5�i�Ɗ���t�R['�
}�%k����{/��R%ԤN�8��*���U����,�1уP�-��.��jm�8j��/yq���lTS��PR�S3��W)��|W'����X�7�8�	e�A�x�v�*��'6���c���%�HTkd�e��"�ԣ�wO6D,m���)&�`�B����i\��!��s�pa��׀��g�xK[�n��/OG)��6>s�u��ώ�,�a�k�O�1�l��=)ӭD�K-��һ�U7������VF��5� cן��� �˷2��-�b�x�'�M-|�h�n�7Dn����/E
D��s�y�qq!�7�i:$��Ux!����M4���L��N�+	ʾb���M(W_�o��1^ѝ=o��L���]gzʀm!�{�6�#�1�T$�]�J�,C{	F�﷣����m��- ��1UH�gF������65Q�GFX��� sZx1#��"&���q���Bwk�F��h�>4C�k�^
��%�[T\6ކd�Fw1���'�^�p�3:7I��Ѷ�:����!�CRc��~�X��v�X!R43�n���K�X�,�E�xV�lT�aҜm@L^��Q
��}�W��V�|뜧��/g�x���?^��n�0�_�̱�I.�0�x��+�Fl����#�	��G(�X?":k��|��Y�Kq�/9]^>��n>�?��f,E��
6�e�)f�G:��C��d�DݬM�7O5�֕� �i1xbO��kF���L����N�ԋkZ[f���p1g�Fi0�YS��Y�Q?�$=4�s�@Ҹ��
-��H���p�W�x#=�e�(�!& o2s�Ň�p���P�Fe��lN W3�����T\6�9�lZ���haHBa�n�~s��/�k��+�*��x�X�Yo&�{ʡ7���	9��z~�Y�;;���5�7 �B3r��xb�.��1�J��E_��������%����,����k�M�tE�����C�_:�[���/jᱱ�Ve)c�|'־G�b܆�(���Jr�T3��m	;�!�d�
�k�[X��UuM�Alu�1.e 5�Ip(CƣW��(���`a�����Y�n�����{V��_�Ԁ}�5>���r�\�Q9���@1��Ó;���GXG���EF���Z��>=;44gA�L�p���r�m%�O�=I��d�� vߧ&�Br$@�6@Ģ˽q�"��"�3�L� �hT�9�w׽M�mӾb����E���[�^��=�/��ȳ�����ć�OF/�6B�t�I6���9S�^��t�vGyv�2���)c��<ʬ�{��G[uٸz�Ib&��j!�ci^�f
�i�}��U��/�G��G�_��byY��o��d2����ݒ{`�_�W��/�jY��K/�t��s��w߃�S� �a��� �h'!������3Qi.��"ƉB��鷟�6��F���{i�u� ]���'���?�E8�����$����ז��X��m�rJ�ᤠk�q�����g�-�W�����~�vLV8Y��9g!5Kc���*y�L�G���Y`�G�ߚV���T�2ߑZ~O��c��EZ�~P���ȫ��(ɏ��������{����Q:��j��������Q�J/"Չ��+|��'���=���n���,�I�!gزUA��/�<hp��c� rU6�T����'qEb%��u�N��G�2�K����U�Q��b�3��fU�ok=BE�
Ǎ��Ϡ����I��>9��ua� �Z>xI-LJ����S߰�\p�y�q j>-�?��z��X͎ D��������,��@=�!��ƽ�f��ʽ ��&d���8���9a�[���L��?��~8�OA�}]~|dX㨪�'�������H����s�~�#t&^u�=s�x-ηU��\g@:�D�6��=�1"����	���|�=�cN���.�$|��]*i���k����*�{���P�����q���>
h����b�-��>�!*����b��h̉����sk��F���*��"���̨�>���hY�? 	��t�9%��3�)Lda(A��I?��0,S7�]��&��;����4�8ϳ�9� �⬽����b+�WُJ�8	3��E����OK` ��rS��WN�Ѹ��!�x���8�AS��3�{T�J�����b:���|7����;������Z�gA�X�JOXf/w����.x�e��A�lͲ�^�����:D���#�-���-P����z@�y����\]�"�/��C���(�������$�/���2�W��u�6�b���K@�dO�g��(���-'���DI4���"��Y'\��P�e�S���X1f�B���h+W������j[w����W��˫A��>�|�[|'#�C������ ���3�?��LL���/s��]C�GT/B1ʫ߼�|�c�/``�AluBKcd�uN��f]��'�(�w�67�f������އ�N��k��G��q��l�_�=B߽���&�FGp@@jg�5jC�`�G�ej&ֱܿ�
H�SUn���M9�X��������&.
L�B!v$XJGZ5W�9�3��
���J~������-�"v�~���p��+�?v��g�D>pԈ1��>�����4����\��%��}-_J*j�
{v��N������$��*$��[�G��y�Pr;}����2bD
�!�{B�ep�����̺	�)�w.Ec-n쉀�!W�"uq��s׀���'�k鍇Je��G�&���H��}v��Ţ+�z��=I�sC�e����g�S_��I*��F��TFI��)~�|{��=�����R{��u:����>Z�C@�N��M�)��Xky�=�+��aB�0����E��	�iȐb.k���meŪ�PSb�U����O�����*���6�Z�X7�Q����l�L,;���-0��S�z��tJ;�3ݗ~�c%)D�%��tV3xԦY�r誘*��҇���TS�sp`�|�����
wLz�	���7.5�fwT_��^��'PFF�m�u���z�I O��vr�t�͞D����>�w����4������å1������C��2s ���;�)-뫡�czO�};�r��W@'V֯R1��4%�ӗ۫r
�1p[?��·_|Ej
�9�����;Ḏ`��u
)����acD�oDժ��t�C�bc��(4�d�!��'�[�@T�X���Q�"�!$�kA�g1�Q@�r�,��aGKA�q<�S@�3��8ߴ���C�,��p�&��fZ�t�@�e4��n�٦�rߨ:�o
@�1b2l�����w��};�g�7@�@\��H�M�9D�׬(eQ�@��щ�%�9�c������9�[`)x�Ҷ2��Z�_6�����H�ۖ�*��J"PJ���1�b���g�u�94@,�N�̕����3��qJ�ͷ�_<N<$$QjeߨثQL;j6N�?�fZ7���\8c��p�9Σ���7��t��
��Bnv�/�U��������ι����_҇�b����	dj������~YQ���;3�	y�����TQ6���qg2�8�b.W�g��8���@�5�n}�U�`_�%��NR���Z�= o���-�D�ఄ��-�X~��K�p�����1c�OU�?�|�*1���I�N�����!.�G-�h���5M]�pi�����1qX#��ϳ�ƾT�:>����Ѱk������65ջ�g״�JJ-\ܧ�C��|�-�8���wn��N����{���K*��5��tj�W|o+����l�WKzJ�ڔ���6�o'�w�8���`S�k�k��kj�U��*�����P|���v����c R��˞R�'�@+'��ZzVD��O�ܛ��.�3���z����1<�g�~h��@�scl��j�K�6�	�\��d��<�ɹ_��_��ND�z�V�!���e����zi9t��h|�Ӄ�#�C1lm�{cB`wj�����F�k9��bz��T�k�8]���f;��/O����?0,:�5L��S�6����ߤs�������y����o��r{4�'1��&T�x��?��f��xE�;M�2u��>���Gq�_d�z��|�Jl�s�L�<>G����M��I(�&��$��*r�T;��5_���t1ۈ23o���ξ�72L�ÎA�}_H5%d����'���z5G��^���J�Ci]-��#��� �OL7�t�<��G[xD��	$x!��o���Ec��U��j�lXa��_t�nwI&#��xLZ��״�5^�n����N9��I�􀛠x\&ꩤ��U㰌�|Yh\�̔/�8��9���`�q;�ə%�,IǢ,<���HE��GVl&�pDy/!��'}�?�VLQd:��V>�gI�ӊh��X$.��3����}��MYc#��S��ݒ���LA��b?�M�B�3݀�m�@�e'&�lK���6*`U�ݱi��꯬�V���ԗU�&Ug ��Sqj˯q��y9?����)8$Q(� �\��4�g�\b���;J� ى8�be$����1���SD����f��"~GJ��i����+�gTZj��8��د=d����u<�Z4�8Y�i�E$Rt�7~�i~P̰�44��sqcM�)�N�����E��B��"�3@A�wsw�Z8�p�S�o�lΤ�Ą'bTSBֆW��j~w{Н�ؒQ��e��̶�����B�x�(����	O+��k`F�&����g�@T�˅HR=�a+�.�5]��)����9H|=ynk�ܱ%��<߃m�&dS�5���9 �Ϫ��D�s�m/�B�g�^����<+d�	�~'�Q1~=�QЇ�@��������4�2�@����H)G�9W�7�ɔ�B�,ɞg��;���� �����[d�o�*�Eh���>{��H�%^�=�!��<8`���Fn�S��<+�7\�\^��`�q}�ʘ&�<�Sw����u���.��15&*��2�@�%�`���9Ai(C�C?��'d�Y��=���-�T�Mh���}Y�v)�sX%��4��Vl�6q�20T,XV���(�B���k��"�A�{V�p�?|{/.�`γ[���1
 < $>�`D�<�`$��v|o(~�O�����p�"oy�IU�Ǽ�2�x�W0��yy���k��-�ne���u'fB�K~�&��v��������������Qd�
�ke���)Ɵ%���}�Q'�O�V��k�L���ު��꣡Ѳ�� [;W^��+l���']���	K�j��eq����M�֚���A��XP�84�nr3�_�m�)m��S�eM�XW7���S���f���m(�k>^g��a��k�R [�t]�D����`���%r�-�b)����@qsV?�a6gCv� r��!=������@w�2���A��b�&��׷�2�x,?�Ւ�wx��_�$ 6E=��k���˧��)ʣ8�+7�A$۪.��_�I����#=���Ų$���XNX��:4B���gY]�ΛFy�&c������OGLO������E�N�ko�.����àB�e��ᯓ���/���E"=nZ�,O��lB�u��!��������R58�-�{���v���[5�Z�d��U}�]o"�i�����W�1[��tV���|��}��t���E�w
����=�nOԋ�5Z.s��/?��NGx�M����S�����F����B�(�����P���M��@5�d�qJ�3�4�1��������w[ZsZ����,�؏�+X7���@��ϙ��VO�w��B���>�.�y+�!>�]�gOE4�te'�Ed+����B�R�^;��sQF�n~՟$y|'��oC$��I+�,��v�) ���<�q�������{�N�-%���wǪ��Ern\�����k���q6_=�zX%�r�_�����;ݾ�B�3���	] 3@A�Ŧ��J�m!A�y>�QA`a��loѭ.��6	�mA������5��l���-�D�,t��'�6c���b\�\��ݨ�
���T8'���4��B�8/�O�H}�e.A����A��ڳ�Zuʊ���w=�Y��� p���_�V��n�s};7�\
��/}%���)�Ar��TQLP�/�UT�6���\W�����8�<�)z�]x�-p����"��E8�V@Ѵ2���ُş�U]~>�>�P�bjQ������������t�HVsػ���Ʉ<x'[�g+�hg�6���"3��0f��A�S&P%r�iD�,ÿy>��	oN��H �����<	,B�^����y,��`���8��'�͟�$qn���ݞ�tNl�ox��|�H�d�3�u�E���ga��,A۝�醌�U�#4���"�&<He+�{-0�=��d����N�Z�yv<ՊM��L���I�_s�ດ����HH��^���!�.�W�w���jƖ��ˤ�I�V`��Y� ��X����鳛�C(g��fz�G�U����/Ýw@+�����X7��&Jl�]�7�J|��+�c�"vв�P���z�1�I��5=��5n�e�8���:�� �se!��yi٪��\<��,厤iN��#\�`d��g���F��e9]��u�:�oA��tj/S(�c2-O�����Q\�miU��Ұ�c6r�TS�*�&�~�f���[m{`��Ì�Љ-/<^y�u�C���t�F���lG�j�"HYU^B_�����o�݈�H<���I�q�2�l. ����X1�sp�Dh������&mae�k�I\T�7Ӫ��X����
n��H<Ҭ�M�������u+y�R��	� ��[��l{	����m�������4q@:�(�y��$q	KH��T�cX�8�t"n_N+���}�J.*��Βd�O��Ar��Z�� �bOWG�!��0D(¡AfJ��B�#�
��榬����Y|k}!��FR^R�I�w�W�r������
R�N*��kK���2T�Q�ѫi�b�Q+u[qSKԂ���.�`*�U? j*�p2�uiGp	o��5[��Y.	����xh���ٯ�B�b��]���V���6�ݍ���
�ϖ�t��c����^�H��1�9���9?渂�X���?~��9���/����s�<6 �M��ʋ<Ƃ#��g���G}~ &��x�&�r:�0s�3���&`��L H:����f^?j[.��^�&`����w���Ǉ����c����:x��x]6��Wu�s;עɋI!�r\꾘ʾW))�$6v�="wi���(�Vr�:�bZJ 2�I��6b�o>���-�=ϊ5�5�� ���}g"!�����]�D�Y����MtFӂ@���UIyNg##5tx\ꍢ*����&���	�MB �+� 8Q&�Z�o��ab���-;2�`0�&<��+uz�WqاX�l7%�ti�����;8/�ُS�}��e:I6	��v��u
0S��ׇ��s^5���8|N���H�87ȧEs����eӋ����!3!õ�#:^�����������������Fq#�ڋ��A6� eo��<�g��[5�znE6iv����G���U1:;N�uk�ȇW1�
�U �LO�Q$��b)�G;s�7��F��r��r4�Ӏİ� lo������(F?
і)��j��:�q4�j��Ea��.�=Sۄ��[B�R���?�=@�(�	�-�o} ۊ�2W�]�sq�J�ޕ���]5�o���ԥU�Ȉ-7_(4�`?C��q ��j��L"�ŉ�������œ�S�q��`,�OLl_zC7;D>r��d��X֚��n��W�|���|�G.����6f#r(?�ѐ5��=m�N��"���o�����e!���V;�����0/6�	��-sp ���HdyWp[�8�׳NIX�_ю�L:Z��>R�o����D2�I͐B��E�|��U�؂�7���}S�Q��;]GD{ACx �Nt���P�J�.�8YB�cԓ�p�p>\A��k_�O�/+��%бlq�U3�ugz������)H����\5�f��yʨҀc�Q9ߵN]g�rt�W(�Q�0l�.������NV?l'~���CT�[?L�,�������p�����ȯ����P6���ཱྀF�uAp��)>�R=��yE:�����$�'th,�`�򐹿��2�JJhʌ%r']!��&��,���V�^�6�r&�'��}��\�*la�\K�~�������U���;Z��X�̏�����u�Y�G�Z�K�ʶ�.�=��><j]��X�pN�[�Wu��P�]#�����|�6QST{ta������k�ڤ+�̮I�)J���@b ^���Ҍ�]���LG�WO�-��o�,ۑ�]���)Kf�V�:	�T7�����Wk���r!��p�Gc� �s���*]%�����q�Z3��7�� ���x$�Gf��J`�4�?��IZyM����	<�-���e�Mw��#[Wބ[>�vQL�3m8#DF�S&݋1�I�w��A��GQ(/�K�SS�YʹI、�V_F�	���H 	�7D"L^T�l��|A��^f�nsJ�Jd,�h I��gjnU`������JAa�Ux�z���"��G�/�ιk4��n����������Ua�RL죴����q��_c9�d�O�ף��V6�t�;{Q�e�{p�k���t�&\���襭���m��e�B���5Ko;q|g��8��H8Y/��*��N�qV��\p)2s�y7��3�Ł��n=�+������3�Nr�X�i5��~�2����#��8Z b���!`w��c��kX+��B��L��rA�?ǿG�
OD	���;�>Br�=?��~%�JRѵ4�|*\��3hr�F?wi��^̀f ���eǨ=v�	�_�j���Z�}������TӬ�����fe��,�����4�k�P�(5@�L):R�����8�Uԑa��]i���M�_�p����q�8�|0�WӺ�b�&t��|�3�K)�H�k�gqVDB�N�{P�t���$�1�H�����)��Uᖦy�j�q�A�����g�O1�ݷ�Wi<~��<^�>����Gj�L̉tv�_$'4��m��:�æ4�_�?�q�dV趨�TW�0�V�n����_=��cĔ=�|��wN��'��LG^a���^�Q��O��@���ut��]O��[�Sj�ơs���`�/3�t�:���!`�v!��-�0pBW,�Ix��&\�1K]����u�����j��f��\\]DY�����?:�6�[�' ��謦�(�8�/��5���?=[�+qwVhR�K
�㡓wuj���~d���NP�z�d�=�3t�Q�M����
��c8��������!$���s��f�ާJ���m��C��4��U���*��c��ȝ�ЕؖE�^'�ۦ�q=K	��z�!lc�5?��� [VO �
53
y�<,1�P�x0�ni,����h�~����e	?U!�le'�?p���G�)4@�/ѨAB�z�嘜��?�]�fj���-JO#�<�a��䲓3|�L�x.4����K �w,�u�!ǂ"Z���"��g���+�x��:Zr����s8"t�^�@n/��h�:���:�mr�/�\���ߑ�CcF���5x7,��Z�dc���|�f��� Ǵ��c���G��s�g2!��,�~�OȀ�ˉ���S��=�+it@r�@��r�'���@Y�Wevề떰�� �2����Ŵ����ڮ�.��&�g�{��o@ZQ_���zF�_�j�&׃�]�I��AF�W��&�8]g4���y�o���2x�q,��h�mB\�#3��K ��doԗ�O���oh~&�ު��i$q4�;5���Ir)h��~o��`�B���/��t��JM�׾_dFj�UrNĶW#zy��͛+���bYr*� �cbτ�ET.ItK�P�=o�N��L6=[�p����6$q�b���y�I�jV�e�<�7[8�6����9���������2
Ԗy��4Ѯ?k3~��$�UE�ߌyk��Yυ}t�r��$o&B{�L_P���@l�u=�`�#[	G!��ɕc`k�����" 4+����
�����oa���~�(�6����!
�t2v�X��s��2�A;,���V��y.1@�H�IX6k=\�U�i.����{9ꝅP���a[�8A!����V�2w}��Z��UݳTևP�F��VMZ�f&�c�j��dڒ�b[�%���6���Nk��M�,�<��:��Cv�Ax���'c���b�L��A�L���7�U�i���� ~�)cE�Σ��2߫Q,�����R:���u�f�d�E��K嬕z���[����ٹ��u�*�#���^�A5ub���KnZH̆�$� ::wJ���X��ZM���KkWr2'9�H�-��	.籬���G�J(8AB�L�r���q��~�8 �2"�y�e3���{����$�����@�>��xR�u��n�2E?[h6x,���r����ciE���>>���1��)f~-��۟O�����Mn�|fҹ��`k��"w�vR��\ܣ��u��=:/;v����j4�(��\3��.�p�=Nr�+�i��vCO��5�显�UV4��~o��#�89P�^��MFuZ���0�ω"Z�A���G���S�n�T�c�����0�!GP6u:X��Ol��,���p�WD��S}��y�<��]���ڙ����;/rbr��_B6~ �@�m]�����e����f�B"���M����q~|~LUN�g�3e�+�"�K���Q4�PY���,��ʌc|*A�c�o�q�؜nN$�7�,�nH��s��#�	�gs�V�K�oiG�EY(cs�>�������@:0�c���m���d~YWV(ӈB޲l \�'���fh_:�8X�p�Ռ�ehO��_�JfhP��3���4����'I }O�L	RnU���,f#l�o�k	ye/�O�P�j�����'9��ߡ�}��|E;�5�Е�\�h���JB��3��ywM��eN��(������Ղ�]Xm<�^E���M�=��g�m{��B�����# �d�\a��N�*��Q;�5�8��5�n��G#9i���lJ_��n�K�g쪄�dJ"�k�@�붹v�q�$;Z�wк���5dֹ��S�U���D��$�Y���c�8W� �����������89�q|4�	�Ƙ?ng��E{���O3pX�_]Gʶˊ6'�`��Tx��f6~��
�kZHE���(��h�Mx�-����a󁝁�cR�4�coy�d)GEH�<�a��!�I�5-�� ��q]y�Ӗ�s�?B�ߟ&[��z+�P��L`.p{��FT�h��cB���:�I���9z�����p�<���J7�8�G	����@w,���篡�ÜYK���)�InA��ʊ�����J-�ݯ�S���:����(�[(Q�ó 6��.Ck[� SI�S{��\�~��5敿1��ýX�Q+xl��pK���ʇ�������n��/�'��DZ����b��PLQa�]D���R<����o�ѥ��M�ik���n���y=����T`�hD�&�gm������x�u��9��)*���`�^��b�k��A��q��Oaz\�a�&{UW��z��f�/�z$�3n�>yP��<wh{���� ����y��!��	�uue0�v�InS�4p��J��v�2iJ䶟���ڔ6��S�=����bt=��Ǝ����.��:��Ι]�Y�m�����P���y��}?�� ܡ1;��G�N.�`;�� HI߽-�\e�,�VG�{�� ۋ� ���_�99ѓ�l�.5-�-P���l�J�Z���z,��&��g*[���L�-A�[N8ԑgn���?��=g1��|q�\V�oކg.����
Qd�M��������˗�i���4�f�E���K4%��Pgx����K�g��7��DVn�L���s��IJ�'�;�X	�H�s�[�XX��Ƥ�E�ؠ���b)��e�VV�[3%ƘW�<�پߡ��d���Y/J�
q.���S?��R�5�;��m'�'��:��p���n�t:��0���Z���y�����m!4�9�]k�i�溧 ]{�#̲�"�xK���L�Bpܒ��5jz�B�Y8X*h�}�@Rr!Y(����`���BW>�Й��V��S���չ��?&�rA�q��f��:����n����	Z������?^h�s��,�](��J+5h�ڋ�s��d��=�u����	PY�5r�����1��n�n� �;p����]�c昚�*45�n�vm�g,)y j>��F�k[��?ӳ���*!5��m6
Z��~��!P<�E@��s������M*!Օ���p&/k�e�[nl���c#��D�V�Sn\�"���Z;����Q�g�t%�搇�;0��� ����A��E����,�^�y��2J��2�6�3B�zb(�}A�q[��������5ǬT�Z@6_QARIW:�����a|�w�׫��5�|3oby�/��aͥI�؞�;\	S"�L��uÖa��TPy�������H��'�R��M�er5o�"C��>/2��a�D���I��=ȸ0��(�h��̻��u߇2����w�uq{d��J�fT�RŲ���^�K�-����1qE
�[<��| �_�2\�S�&��ud��B��P7�#��,0Y�GlkV%�]�q� ��Z8�P����>���]�Fky��ACp��ɞ� )�S?M���V�Aۦ!��P�P|���[K�Չa��T:G��B�q�!,/�,�fM[�ɓ��;h��JcM���_�d1x�-A���W;O�6��Jv~N͈.M�-��ßدfߥq2u�3�<���;�j���@��t�+T`$A���k��K��d�P��x606��8)5e�FV�F�t�|G�&3��y ����?ʺ|C���4�x��)���ж�K\�(���<�,J�Xw�t���?�h���uA�X�4{	&[`.�H����r�(������z��lU��	�7]5-?��{-��0�^��)�#U�s6��{U���=�yHQ.�9�X�W�ʩ���YR�\��29XI�	�D�a�⽊�&���c��)ɇN���l榧�y��=b�YB�-�k�q������<�@)�<2�tSh{(SS#���.gx�S��#�����B0�.�4���!�g�6����<�O��w�<jNZ1h�8����"j��"�m���9-�����ؚ�эdp\C��^�<�ߕ�G�B��Xڽ�"�k @FQU�T�=o��;+�Ü�j̊Ӗ*���*��w������2摉t����Z����Jc�f6n��J���J��L�O��N3rI�U\$��'ȽG���t@'p(�!?_'��WYH �+C�l#�,7��|x?ݑ5?U�m��	lf�:�^r���D���8�t�a�E�$."5n�U��n��j����ף�+m�]�;�������X��~K}�`KwQ�_P��\��ʓ�\̹���	����ԇ,�� ��ed�QN�9�;�؛ʧ��~��Fy��3��D�Ov�@`����$�����{ï���I%�A���Ǭ�-i��O+����9F���J�˃�$Wj��ci�we1�t*&�c$8/5��M��!��O��=m� *e���D�e`y���ʤ�_ؤ ��#�`5�.P�}<#��g�@�gu^�_������:8��7���j`&f���Z�2�Цh
�W߭H2��/� ����ҕVR?���G5�Qք��t6���p�7g}ɪ��VǦ��뭮��)�_g6N×F`�	��*��?c͎�zx>�bA�uٿ_�J��α�H$JH.� q�jxtfk(!�w���y�pHs*��q�-"�$!R0���yt��ڈ���!��L��n�6 �_��-����� �l��}sy��D{_$���%������fE��P�l�Q70��<K3��L��a"�s�˾�Z���4�D��>�~���o��l�Q���,	jx��S𢩥!#�k�����m u��2�q��a�Z�zD��2I����tK�B��P$rL�b�m�`Y7����E,��K�]=v���ǻ�/�l�	�������[�1��MFnW���@����e��we[�?>�x@���`���G�,�]���v;�>/M|�kH�d�Cu�/�
�ǲ�����*�ݛ�m������jO`V�����y�O�� ��*5�d���~�i	���O@',6��k����_�2L�(Rp������[����ap�l�	IZ��ށ��O�ǅ��?7���
b�=?f�C���N��N���Α�
e��H��T/��@��6�,�悧�ܻ5/��2]lC�L�6ΰ��)����Q�D���� &���Qd ��W�z8�6ZO���p�����tX2��p6�s��s�����Y$_��Nny-52��2��Ia)�3��i�>W�h��/��%���4
��"��ޣ���
��pثY5����9k����;� k�c"s�0Ѥ����Ki�����x�Jq$���O�r�?�Oj1�A.�Z�N��?�����t��K�T�u�ެ$���*��o�!Ԃ�5����n 'cXi"��x��'�[W"��ۿ��wUt�&��q�Q�τ�K2-�"�ӈ >,�I(�9�<�e�hB�ZE>�ZT˛��S��HT6܉;��@զG���V\�������ikR�^MǮ�&�n-��`�5���#�5��TV	!2����a*�Û+�5xz�֧#q�G��v=�;�0]��e���?� ��f���r����e�?���
�q��Ƀ�0E��gW��=7>�;�����BW@b�3:���I���%�n��C4���mőuu��2XboC9C�O d;rx5��,������Ĭ�D�[5"(�(���3��[���B*�2��f&5��s�=z�Hw=��W���g�x�Lğk����M�xB�*@���K� r2 ��2&_'jrD�l��B�)�ii�/����[�8��*����~&���H�.:/�eF��.��1��ǉ;WڸtUt�a��5�,��jK��uR���g� �ǑG�1������r�����������.����_���E	`,a[�٩����aA4f���Lن�ԄO_:�X5�۾�^%|8a;yz&��P���A-��n\�}��;P�ה�
�j%5�Wg�0-���b!T�:0�2���u�_#�a��S=���)(�����yp���Y�^�_��Z9��t��c��e���xw��turD����E�W��E,��_�	�0vI^����Q{o�j�?8=�oC�<����,��?ز+���1^�:�r�8��ņ��b$5\L���O|K��=2�f�f3�f5uR��I��8��#��q�ˬz��	Uwm���,�Y?�����֔��k�-[T��x�l���y΃�W��Ѷ��V���	�9�v���3��f�WȄ���A����<8dw�{�;���9P�3���!��&]0F���\�����n�2�r������r莇CP�UnO?d�*Les���]ж�y�	�QOQD��Yb�h2��a�~��ũ�{;�6�#�آd^	�[����_�A��74�8P-P���>���Ӵ�Z��J�K�bˮ�սy
�+0��J_(��7x����,(3}��_�,�&�܂�[,8V��!J��e�f96��ˀHg���a�*�o?�@�͖�Y���&�ˁ�s(�{d�'Π)���P�����'�7+m�,�5s$���8QUF���qɨ�J����Dʅxu▧y�(����vD2��A�;��D�A0
R�Y�^��$�71J2 �C���j��ٙDy^��b~r�Y
�����dP��h���Y
