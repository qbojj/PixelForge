��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0C�V�D㰬�hBW�b�{w~�T����#�e��Wb樘!zi�ߋW"�m���)��ĘI����Z5M��y_��sPi\�M��HG�6`������/���S�A��n�Û��с(^���.�JN?^��h��/?�Z�x'4t� �V��7����9���I7�d�x9u��� ~&<�?mSDyԦ�ġ��:)�����ǰ7?�[֊x�mnM��xڻ�S�V�pF�R�zl�XC}�y�l�]Ƴ�"����K�^r2{���$#S��Ȟ�Jk��G����<�T�Kl���)���&x��wW��k���C���0�F�� �F�6%��(�l$��J�U���U9-�R���;x�.X:)�%�\kB+�c�K����4�Ζ7���
R0e�<s�29�S㻬��0���wG�$B4���0�1��Re����t��zg$.W��)�xV�\8+������ܮ���m�Z)W��S��	|�&e�{��E�Eyd���Xy��m��©6��b3j(xfF?.�����`��E��2��[�59����c�Dy��MI?�b�`��W�4P�Ŋ��SFmPI+�A|w�(.�1#�1��)DF��뢪zI�u�y1qw|w1N����,H���C�����!���pu�2$�./�^Ǣ��K��6V�no�v٦ˏN�\�1���B�����H���t�V���i����]�Y�/�~�;�k�(���!$�	�p��
h��u
�4�]UD �b�� ��8A*�����2���"V����fQD�[	X��6ܼ�+6���3��
Omwa�k�� @�����|��	bYGR���Hn�w�)8�@�hds�J7r�0��-���Ҝ����h�_"l��(+�n3�l<������]��]�zA��j��Ԛ"=)rn��M�%~�lWG������ؒ����vP�M�W_��P��}��O(����~��  ��)zXq�����p��� ��ʥ,#��S�~.�YGkK?NƇ�-�L(�(����0Q,ɏ�a=���Lý4�ꘘ�ʺ�˘�|��5��C��;�ݸ9A�&/O��6/m� F(6���
Cs�^�)]����T2;���0�|�aE���3�
�+�V�O㋼ ����5Iw}jq��S��Sk�ۓ�`�Fρ�_�J%�A���p�"u�{8�J�R��X+vBѐ�����Z/P�Q3��C�!��E~t���^ޓ�\��?%���-T����S�L�..d��B��-��8Ө�p�.v���<m��; ���RF���^��(>���{6xay�FVH)��^�f:�Q��k�H�a>�L������ �HS�c0��������OL2\^����Yǎ�f8c�z�f�������3����(�Ҟ�\���*J'l07���k�D�y���#;l���+]���C��Uy�y�h>Kml��Mrz@���>V����I�P�o�H�ٲ���Eg��2�k�1�m� ��N�ŵУ?>����?V~�,�$��C�!���X'�����}�'H�'�a+��ێeC!�2J��ф�e��	:�}O�AA�s ���K�ė�c�q���օ�l�M�K�._=g�
ԩ�'�^ue����]��7�z�N��ϖĲ���8��sK9�n� � �[�U�wY'��w��
!�y���|�텙��be'�j�ү�����	��ӻ¥p�b0ﯷlC%\�v{��7�x����[��6���4���,��[��g���䒑�j	ƥjVb�4Q��r��=���rn�98 �o�D��/l�*!��n��.8<8ܴP�_�nx>|��������`�9��k��'/;c
�M
��Aߵg�AHU������q�}�_*hh.y�iT$5����s��$԰I$3|g�OAi�<\4y߄R/��iN��WB�ضѫo�*�ם����X[�K퍬��l�Wk�\"�^kü�_ ��S�ig�Qz��T����*�������!��qsJ�K���6�M����q��ҙ�h�H�
�\�k+�t[�"�9�d��5\�E�*]O}�<�=A���:����	�`�=���~`]�wh�#jmQ9�q�jv;�����D���Y���;94r��QLqȩ�%�TE ��wJ�7�����R��ޏ�4��}�����������z�A���TWc&{^i4xU�z�E��~��|�]<zTyQn�3��N���c^���M/���CIzNF���~�(a��!��z=p)[��N���B�;�&�Kw|���ue+4zc5�.F����Jx��b���	&�ݡ-b���Y��S(��T⋯[���,����E��)�|�gn�x��ܜa@(k��!!a$z"Fl�ڇ��-V�����tE<u	�*��G>ɛ͇�#C��ޭMK5�V"���S�h*���_�#��j�j֓	>w͵����}�ZB�~�B����DD��Ol��9�]�%6�vw%�#��lOj������hq�N�<x  ��x�4�ge�j�[RӼ��)�ƴe����Ic����Xug����'U;EҞu�g���5��*�H^�<g�������D
5bK����R�-���ː�%v_����Dߜ�}���ƒ^Q�&����C��	u*b�X��3�?��B��bLHЛk��&��d�84��K��Laڌw��1�0�ZьEקh)��.��P����C�i��Q�bGw��&�x�QAmlo9q��#�z�v>3\��ln��[��z{.��.�
G�+�(�&o��Y^�u���2�,�,�%c� |ҩ]�a�ߌsa��aL��zh
��u����o:��x�׳Z~�Gɛw
%-T��O
fFh�Do�LN9Ը�݉��@��ܟ�^��+�.�T�|�h(�WaS}�D�&���{e��44������)@VL1��1�D��$$HP�:^]�.;~��Ϋ�Y�ū�Q�Y��N�E?�$W@�ǀS~i{�H96[�6B�t�Y�b��UB���T�?�=���	Fd`YC�S�)fHq�
���	���E�Rz�����l�b|H	l����>�j�x�k?}oW=s�w\~E+˭ m�M�^����^V��a�0r�*c�&�6����ݨ��	��Ԩ�L:��D�:���Td�?A�J����i�$���K�Q��M���!�i�#D ���&����V!=�^!xֳ�r"l�G��WU��}�,��S^{[��#�#��	�*"`�*�!P�z�2�ʱ�ۭ)q�v����� �FũAK��_U�N �|(�&h/�iH�LauD�^��-;�e�<	���/v�$m1D��w�|�ԉ9}�4��W7�:�~bQ����p!�L���]�4A��R�
�Jˆ�<zj�+����<U@�5�����B�� �:�)��灆�{_���9$��e�RE������u�Z?W>�& ����p�8�+dX��ć����%��d���ُZ�gn٣�d�I��y5���_�&J��Z�������Qq�􀦲�2�^�RTD�3�䞙6c�Ȯp����Eܓ۞�`P=f��`2h�ނ���Jnޏ]T��e���=�&�k����'Zױj��+��f=�`tp9��O�v�u�����O,e��7��F5���iԼ��	�)gnT$����츨Br/s0�k��o��c�_��Ue��c�Qv��v,����'ek�������iV��%�%<-8��7.����P�����?�W�	AN|`{N�<Ί���d��F9O�	E¸!��\�I5�L�9�����p��Rfy���=Z�St�%��T]��r��\lOsۚ_( m�7��t���zX؃�
EA�p��d��dM��|A���(�:;phQ� }2�C���*�#�G�\�V��x6��[T)L� a�ҙ�d?�$�S��u���w�٥���ߞd6��/�n��3Ϧ������78���P�"rMt椅�R��� ��7�l�@h�t��/ũX���\�a�S�U!�?�12ѣ$w��VX��;�Cw[�k�V�߿�{�V�i:QqQ:�t�"*6&D�u
2�T�d�^��՘�<y�Cƴ�_=�4�9�Ǝ"�r\��{�x�,�$�P'�=&¸hɆ����ިGIsB�Wv�Y�	t���l}�EȦ�Ou�]�]���'�.X�bQZcm�Sm�����7"
���S�X���Us���w��"�LQ�32��1���5Ƣ�,��Ș�o7�@�X���(AQ��"Y�H�8�&�rƇG��bC��V�����p=�� ����2
WȠ�hǅ=�~/!����[�N�t�ண^Ф����[����U.Z��P.�����+^� ���6�Ѿy��la�k�'ro>��^��OBU��%ޥ�D������&���@�����ل
���фo�v���W���i�Ӫ�FW��=�~����$B	�`f�?M���S��GwG�m��]Rѱ�6�\و���/b�o�]���j��3��f6���2���܄Ic�1��K�����î�B�����:��P�m����G�2��+7�{ns��1�Au��~ޒ{댴��̍%E��	`�����.W�^���=����o&e!_�d,����k�ǒ�����N���{�]E)�0�-L��t�*l�(-pU�����m��T���!	3bj�t{-g�-����◡窿������� %l;�lS�{�r�(G�D�K'�Ԉ�	e�OZ:cՎ��d�,xM�hwk`�\4[U�����wİupٕ:[��B�͞{�l�<�o�
���9����t�2����t�Gz�'4��v*O�Gg��J8�����(\�8���n���Qg|�ʣT�_��^b�h�Q�4�@�1����V�'�u�ixtj�Yz�GY�;��6P�h�0<4(ذ�?�h>�Z��\`K<���|�]�Or���F�|��4Lڛ������m��]4Q�¶
��H�8q����Q'W
�Qn�T�j����8�Q�D����t
I4m)��F��'E��V� �A|�^�^zN�B$�q>�+�k�����+6D�*tx�G�.�MY��H��?�r�?Z���A�sϺ<��O"�l.�� �ŕ��l���*;ض�'��SwF7l��)���FW�G��?�W���T� 5���I�C��gl`�ܻ�u3[���j�k(v�c��UL��I8�ޕ��E�C%p;m��9�\_{w�ֵ�Q&6H��hZ�Es����MvF+XX��?����
�`����M�&,��H������e������-֤���W�r�wR�Z ���ڏ����[P�i�k����`�x`~`�^���u`Z���
�э@��F��iI�bQ��lQ����hª� 'j<5b��.tr������|�D�+>i&�/]j��!{kt�ڼe쬹����C]���*M�шH0��4�����.�n$�۷�F{��W�ݺ��ߋ��22�kW\��4��jbqDnL�?n�,!` S��j%�F�ÀW�Z�O05A=�$�kVLkž����'bX�h��;�6��b����W��Uit�з=֠)�PL�lG�c2}N#�%�r�r���?��,<��E��-௲h�e�1�>.�=�9"��e�@���P�=�J<�n�(�����B��rI��q�������XZż*S��_��K�Dx��~wA��o�@�����k|��[�[�귶��=(V�JXo���R;�>)c�A�9����ͽ��G�瑮 �2H���E�����H���j�7������-�8OM���|�.|E}�e����<�0�G�?mG��撲��d���8�#�����#�ꁞ4�����tM�n�����BUVtO��cٲ�ǜ�7;�������*Y��v66D����-7emM�xg������Q]�9�@s���k«$!5���2��v.`ժ</���vO%'�QjWc߄-S�"�ɷuY�I2N�����8\_�˘�p�@Ia_�PI�K�&:���l�y�+JqmJ�悥�����,^���bW�C��ޥ8���L��p&���yĴ�Z~dDj� �픭�g�RlS]�(j⚃)Y(I�s����y�	�)��SԆi<�xPΊ�S"d�U�����i@�oӸf��k}t��#U@�'���}����{�RLr�\�����y�YTdt�6�pP���]���?�w��]A�q�*���A^?0���lD�£@m]�$'�T����0�:?AKF�2O_�hᚣ�P�?L��y�*O���g@���D��.�%m�g4������܁-�m��vx�:!���M�d�*�'��@6�uY���_�+H��u�=�(I��Ӈ���]��G,�w>P�u�l�}HRk�(H8L�-�=�g)Dy�f�B;~�TX�I_��<�6êţ�k�4w\6Q���-�1�ۺ����Э�U6��L�wˋ/�ɝg�29Wʦ�/Pj>^3=�s#N��ʻ�p�&�Im�lz#���<���6�BS@�|0��B�:Z�4U6.�gv���k��R���>*�2m�G��H9���0�D�hG�^����g�h���gJ�W t����.�I��_�N�F�����R��(.�p(� �@���bZ𑄃\-�&��xg�����=� � ��ʆ��A��#s)M\��.��w����U�v�ơ}�s�kO�(���{��	&�Y^�T�ڿ}��J�\���HT}���v:���˧p�]��ޘ�$8���"�G?������ȝiƎ�s[MI�)�&<	r��̚@�a9���������G$��R6<�k螔\��խ�]�o��l�̦�E��kH
Zʟ�o�7�����q@�,���	ӝ�j�Qb8r��2s�S�y��gc+�y�_��Ӻ��z���ƮGZ3��9������A���C;����]�&�8Ӻl�q��f%�h�����Lݯ��)�L��^X)�&�$��EU2���~b�c~�B϶��'�ƺJP[2�����q�?�(���h3?C����4��Yj�c��x���'3��8ƼfQ|�9���)��W����U�4dne�����IO4n�ǁ������8D��qX��|۬V�2����٦�]��+q)��)�Zy��Nd�cWM�엛�~?���+�@�I��+����ڒ��S���9V���B&I�>�7"]s�~M�T��3�'�����s��:*$������k(p5�r1|�<�����'�a3G�~N��a�K��뚧���~�O5����A��`�)Հ��P����'A��I�Q6%��Ӝ�ƾRA/����Y:��m-:-K>�EB 䳱�01
��,tu�0����J�L�2IlЈ�__�h���3�D��3 t>���F�	���
kxC<K�DIMSߺ�[	�SM�LNv�$����%����G��͗
𷻊���cW��z��Zb]v�d6�؛%kR��=���N�*�^ ��q�3��jn�
��f�d��I[o,�9J��"W �~�p�Cr���7���P�B��N�}�h�B9oW7�h�	�:)E��Q�~��������a��ܮ(��rދ��-� ���j�X4����̑rj�{e*6��*�������4��̂�Ũ�=s�ڹ����(m�ÿ��E˺��%?2���G8{�3���Ι:���ʠ��A�@7�r�������+��(��y5�)��o��C���� ]�T7��j�� L�dj��X�KH�Kqbź���dM�Ho��=�kq�e(��(�[ ��X����=��l[�֭���{0v?����X�ݲ�_���)$ҩ#�Ќ;�BQ1�.�9GM��-�ox�z��'��I/�����K���G3�c�ĘH������ҍz�%e��Y�c��ٗ9�#�S<3����Ϥy���"�YdlQs�>/3iuxA�1V��!�J�qȅ�L-߶O���*h�+���c$IRŻbbRwd! &��Xґ��z��Ue�N�$Zf*U3��!=�oxB_��DaA�혀����������ǲ��,��7���u���q�[D_�(�ѷʲv)`���Q�7!?��#D5\r�~��pS�����F�zE���1*�涳ոG�m�Ͼ�2��s��Z�W��e��p�+)_�����U{�>�t�Q�(L�_��0��t��e)���3�Ⅽ1]����q�T�7��2;����#�@5BD�[�w.(9!p�M%�������h�>[���YQ� ��A}�2�������9j��Ä>6��g3R \�zϏ~��v���:,�Mc�����R;,�T�4�,	׈
 ���Ҥ�~Lp6�J��"%F8j�+z�%)c�"�v�n���=�=� <E���g5	�uҺ��;Q� ^z���- �ڄrR_n�G~.��g4y��
�\j��yBx)*���j9tW+���b�W	���{(�$�~��⻍�{��N4L�����_�Q�
7��[��'��"�[@�f��N��\�db��:��ꣵ֬n�R��	����v�I$e)Ln���r;
���w�ޤ�p7�.WƳF�Uæ^O�V����%��Ʀ�6�8�v+���)f��y��YK�y��CZ�`��7&x�:��0<C�6R2x��D�!@��ONM�샹��ГM�!���k�Ξ�����h�˼���Ȯ�)��):@���o�:�D�v���(ntR�.�\�!Y�tE+���*�q�?6���24��'b�h̵�OwX6r����3�0ˀ7b�V�j~�,�ҥj�¡vO�����oب��b�Grc�U��mҔ�|��W0&$�?T=e	-�&��H�ao��0��d��b����;r£��T�`�|�� ��z�=���-]�?$NFuY����uŘ?��#�=�;��rG�p��T�Bz�;GI|��dˋ�E�" �G�|���P��͡MtX$�3�^�N{��W�&�]����� rE��KrX��8���Ҷp?o���-���'Hm����ΏJ��虩��]/j�b%`Q��F^�O��oO�b���?s\�%�Y����s�����o,�������o2��MA�\�C����U�/�՚�,N���!U�dp�K���T�~PZ<P����T�_��l@X��/U2�p�xHX ��R��#?������a^�#S|-��o�GqH�Lvܳp-WS�k�dN��!�nK��E��~�&u��?W�V9�;#�M�*�?��,Y�a�̕.�����h��±�|��ȥc��ג�>��Aw� ��y���,�ǣ�b�Cv�v��L*P�}�ꐨ�;�ǧ��+�����ht
��A7��g5&Ƌ��NV=�Qų1w�yt� /d�7���I� BS�K��oF��L��r1�:-��r����g|ڷ���S�'�W�l�?��;A�{�F�Q~.go4�E�#��&�yc�X�l�t��e��w'�$�{zf��3���sF7�o�����W�s�����r����чa�և�[��.N��l42�8�%��{T�!l���l/�i�k|�A�1
)�i"�@��2�0����4V�g��u�$as�����{���c��]v�;V��,u��DJ��-r P%#E��)]zZ�Y�
��k�Ո
}2�|�iӏAn���ĕ,�s��.�{V>���m�؊����O�.�Fk>��O�H|�b�{Q �Hq�U(��&�Z/�&p`_��b��6:�M��~�!�%��I8��jS�d2�����5�ެ��,L��B�T��צ
i]h�_z�ۨN!���6/p�%��Z��r��/^m?8��_���#s�Yѫ^L0���u�p����4]w�0# ~r�T��Ur�G�Jn�a_M�~�� �L��0�6��q(�]��k����\��i�^=�� z2���E
���������ɑBݝ'J�+� �������)�p�F���D��M� ��փ���ʎ(��=�R�ߖ���Z�z��c���ؐ��D���|����n�Ӏ�GA�jԀ�﹪k`5Ώ"E���z-'{��;S�{j"�Z%n��u�^�+��$C��ݷc�j�����kyWF�[���!"�隁+��k����;���n��������xO�	酵*6��T6Z�����Z���X%���R_�.�7{
Ї���x���[��F����4>��y�#���]���, d��
���eI:�>�M頨ޮX �fK�C�P�LQ#�C��|퍚���\Y��J�����b�:���m9������^�[������A�!��[l�u�����k����:�a0�Cts�̋GPfc��-^�+q��-�����[Xa�R����d�GQ������L��E=�����B2U�Iȼ��n?k�ӑ�qzVd�ޡ<��'��0��~�H���-a��}�ޗz{���������q�r���b72�,��n�d=Cr��܀��)tJy�Vg.W[`�.����12?�b�
��vV�0�c��Y3���4
g�}�q�:��C~Ɓ5(\�9�Klir�Ħ⒈��\��rO��������� �c�`rg~e���#�_��v��+�P��`Hs��e�H��Np���ܩ�;��6ݍ�P��4��#?�,ܼ�?�'zq��i�]�I��A9���<� �I�h��M��f
§;�A$΂@�n9�U8����ܵ�Lz}V� l=��u�s�����Q�c3��Ŷ�7���@��k6*�t��<�O�]<T��S�!m���l�'�ݸ5�Y�Ƒ'�̱7�����aj໪t��}M�i�aL��+:ܰw�i8��q���K��@̻�>���_B��<�mu�Rߙf�f-tx��ϯ;�J�h�}U�/~bw��c�C��X�ӂ��'���l��slݭ1I;k��Ńd���S �>
,�
+-�R�#2h��0�8��W�=�ԍ�Y�[�����k��[�ʵ��q�ӆI�X�����1+�uoRTkŃ3+́h�giVWH�g��,��`��m�]��,q�,�Vř��FC�A��\���o�GI����<6�Tڞ�<hT4�J��p�;���2a�/��Y~V�ޢS�lG�%��*|a�h0D����<(��$�Ĵ�e��]^��`Ri�iJ���}�"[�(ݑrs��\���������Kr�e��@�cȒb��m .ŵoN��h���.��:�7=��!�Y c��qW
��ً��_9�An��(��������Ɠ�ޑ�� V`E~2���I�)
�p�����OR��:����yۄ^܎5�Cz���i��gt��_�#��Da��m��qV��*�.���t��;Ż�V�<1 ����x�y�h�Dh4�5^Cz����!��4)��M�W����ծ���+�X^5��W�.�ATO��N�Q��:�I���.�z!�4ج��'%�JN�#�ң�w���E	�����(��#/UU�h�TPu��K���nrĺ��&�̚���ؿ���s��`Drm��2�/����R���=�Ӷ�-ax+ӵ�)~v�<�xT���1�����E�W��^���-2�G)Jo|�E,���`Fm:TҼ�r��[G*�Ӑ��نp���T��o�1�Y������:��>�w�����rT�nO��etr���Á���74�����zǰbԃ�S�Ǔn���"Hx�|�Bbڡ�Rtzܸ��G�Ob$�n|☜��r��}��.��鰜�(B0[9�r`(�_��7g�����ǯ�`rIƢ9͐~�ա��W�����Lu�y��������ϳ_��Y^y�k�����̾y��6l�)[��OC:+r�,���$9O�ý7��=�PQ*�q�`ֶ"E���P��+�����.�!�"���@4�C��U�zHn�p_���-�Ο�߮����(o�@�n�K0��&�6�H>P�l�N1xg����:k�	^���
N?��6�<�Po�װ�����خO����9�;�o�� �;���8"�B��4���������h��MBV�Ti`����|u��}�����R�h%p"�4�eC�+��$�PG=E��KF�*�/�s�W�����S'k�2z��П�1α�v�ֲ����fy�Ŧ��!���,{z�r��v���� ��m�ZB��	L�m�.ђ���O���M����Us������7��AՒ���^:wؓ4�N�
\��j�m`%�j+�C�r��t�Ho���
�((͏O�ЂIׅ��{ٹy�0���T�
����W/c���o�6���6!��?�5��k�b��K�X��,�dk��]a�h���^�Dpn�F��%���z�����֑���06ч%����4o;�Ht�΢�>s��'	�
�@�~k�ckP�����Z�"ޑ���:�	~.z���h�B��F�>󴕢6�`���ԼWe�������9�> U�Q�e�U���=�q�$�Nm��R�Z<��f���[�C<r;��`ܤN������s��.�؅��R�)�>W�.`�|���u���a����\p*n(3�
��$���;J���wg���0&�r����Jou��S)�;|��Ґ�=)z������:vw��p�ƺ�X~ھCO�y�ݕ��,v4[�>e��"��G�)��h/V>��� <<��0�a���l#���¢��e�Q{�K20�$�B ���/����¸x�k���\�73� JWfx�]���Id��A��T9�%XG��/��2�!%���ꎁ�seS��d������Z3�j�۟B�t ��d���m{���P�@��4�'
����,��r���CVl�ig�E⪣o��3�C�m騿�%�Zj���3z��sWѨ�Cq�+,R7��!ŭ�Pud/6W@*r o��Z�!$�3-��f�Y�uhhT��m[�K��1�'�_�DW��MQ�|�Kʾ|׬�����Q�a�d�������vwq�mZ��LOjzέ��P����
��� _(��]�_*�ehnH�� GuT����F'[��[r,��N�7���;q/"Jrt�n\q�}��^>�dL�.y9r�Ѵ]������K�/�_�ܵ��]�5����9���!�r"�ᡘ��&��A{�0�m;���@�[LW+9!N�z6a������r&b��tR�~�4B�I(��Ǻ�#���L"�-�;��-8���:>}	r��w�Ϣ����3��7w�۾�|n�����5��x�X�D�~�z����҅iPOu��Ʊ_��T�g~Eq	���w��K���L����A�Ad1�W~�mI�2�3?����r�h���(��Izu����cvM4�}��Ț'�FU,{(cK�!+�GI�gAL�P������ҍ��gv��3�qV]�e�<����U:w f��=�Aۥ0t�<Q��%Փ��#O�U�.�� ��X8���p�����V���WV���P�Qsvw 0�R#��|S�&�r��l>F��t6��6��Q�/HC9tê	:���*n�Q�?e%�&��������-���6`z*�A�1���G~D�����Җ'���������q�w��R�H��*V0;���2(/�Jݱw�F���>�o���=�<��+?s��>`���= 9s��'Y�����
,G��58�FS���w��9K�W_�S�L�X�BO�� ��ѭ�|�ݘ��j&!���vLE������낽�y[)���f���� )���9�ju��wޣ�v��S���v�5����?���/��.[�w��6�D,-�ưZ5��M�j��7�#�r�%)C܊��Ԕ�����[���^	�Kr�'�J��t(J�jd�L	ܣ顐�Ǒ�F�"[G���!=�t��;���JkI�j��td] �:ʔ�Z�R�eÂ�]Ot�8"��H��ЂLL���AO��'P���+�/�0ef�*���������X,5.��7�'��E�Ӱ�Oc#JsO�	�;h����e�s��E����!��e]���rl�R��,�\�	)qѽ|(�)�A�6�ZE���(�s��͂ �ޖ,,�n/�J��.��M&�vb�l/j���'8_�R�����W���6���b���N���(�����5<Ǉ2(�� �	���T8�� w�ݥ:����U6%��N髛E �8����}.r@�t����o�ţ����JZ����Yp~yH� o��釀��-�=��V+2���Qa&��{�Ŷ:���Ȗ89Xahb���Ҝ]�hj�GN�������.�*t�U�����qt���&T��|<�5����<V��em]MTvRF7�U\�Ӱ)r|5@��t���o��2�͉zr�u�1�-���ڸ� m1�`��y��K�E��%���4ΕT� l?�W��k�ȴh�<�oM>4H�	���N�q�'��o�h��|c�����k	�T�^C�?i#axҚ�Hiz�B؞g�Y~PQ�th�ew�� ���?�)~��Ѡ��z&�0�Ǯ��œ0�NFlN-0�D+D!Z��C�>n8�ihN7{�t����O,K���2�P)�� ���`����Հ��������w4�T�C�-Y�g����2�F�{�~9+��7�	�I��������JΊ���/@���A���K�N�3�9B�d��F�����ޏ�vU��L㯃��V�C�?
�� �� �C�=�rS�%���(?[���)�Wӽ�l�^V�m�pcֶb��d��'�q���__u+���m�[
��l�br@`�e@�y㺀=�G>�z@?�����#����[eZ% ŝ�}^˟��QE�`��!��S�ٓ��VDNF樟Y�߬�5c�}=��{��e���ē��;����/rC��?����=�EcC39�����(��(W�eu�����ڙ�d������׳~�JL�_K�K8m��-� Wd�K�H=�z<H�9b�r�?�o����GWX��=W�lIe)K�i�%����L4��!�R ~���h���r�- �@�>��>_߸Ư~�ID�0���GO�l�Y���Ma��i��؍AїX��R���?��w��Vv��]Y�҆G�ҟ�z�Q�������pj���b���#�]s�sx�G����5�N��f�`���"in�y���ڛ�GF���sd��&�o�̻��*��d�T"����^S�F3!Rb�R��l�h{��,���N�h�i��	��_~͒(�:x%�*����fdޕ��L���1���V�����'J���Qc
��r}�������O��2��.����b���&�_�&o����£�@�_��������O#���ީH�?��RX�x��?�%����$��]: 3;�1*�)M!`#a;��J�����&/��9�9a�¢,����__�K\���|gom�������<2Hl5@��þ��W�q�y�M�`���M~�d�L|�����|��d���<W��;����Qu���5���.`R��(��GQ�Ru˴F�IɅ���H"Q�������V�t�w�3R:c��{֐y�:+����~2Rl]��y��O'I�ۢf#�?e��駺�������*VZ����B��`P#����^�����ƃ��[��C�搻M�� 9�<��#6�=�>������e<b�n�B�(��z��{y�O�w�Zf�p�LhG�ގ���r��kܝ%�p�C�x%�SL���,J�a!C�R�w�},�iv&q#Y)Y&L���L���J�B_#��f���4��@�L"��f{}������n��+>�]��:q�*��(��z%|y~�ހ҈0R��b��w>�d� щ�	ڶ�-�k�~��V@����f���-J�q��q	�	:4v��m�-փz3�{�遝��]�*��c��r8q��T����#��OR��/t��y�\�I��^���4�HM�/��e��VR�S��
/Fo"0�Ö�����9���[��� z�Ӡ�k�^��h��L1= ���Wε�Ik�RiK*bV����rv,Ǣ���
�����$1(�4�?J��O}X���p��zI(?D!ĒC�H��ғ��N�/�ꢹԮ�R�vԒ�ܼwȩ���.sD<F�x$�����^
�˚��p�Vp�>�J�������O��/790_��Q�7l2������0��Heưu��a~�h�t73�[ʴ�(�̙⊃�nQ��_�
�����O%�웣)����d��'��7C37�{Qu��c_e����T��v���t]C�v��[�;?���Wh�;��$�V�U�G��8O��W3�	|��Q�V�ƟLe,�gRe��<�(�C#�:d+W��R]�bR�����lǾ������j8%�8�	B����^���7!�N?3}g�?���w����5d�����k�����	Y�w=��f��Ũ%����|��;�B����tX�6%T`��bݞ�9���� f�Lv���e��?�5�sʷNǝ�0�Ϥѽ����{�v;5�&�y�� 8ȹD�D���@<�*<a*����:
�G��C�n�R8F9{��� ��d��w���ِ�s�m��n^���sy�~%T�E��泥>�<��r��-`�MmVe]x��}!84�]��Zy`@eᇃ鷒�����T�U���/��;{������j9$��8��5����U�>�	�t�L�X��wE&��ꎡ����*���2��V�5�x�S�ۙ�w����%P�F��͊�C`�f���Z����/\�Չ��3�&�ey��r��謖s��wR�8��OU[��z�'뿸��m�U T�uu�NUxe~D5�2S�8I��i[�n��bg�A֋-�ԑB����m��#�a��0�e#>� R^t�	+�=��b����� �-�`��y�#n��j�mr����*|�)܆8U_�:\r�C�T��4ш5����H�"B���� ~H�/~:1����5B�j0. �C�����oT�����j%��?/ԍ���]����(����eH_��ۉ#t�Z-��wFp�"a$�ʴ٫��Y�;q�X�>,^@xv�aRk�I(���G:��9��Pvb0�Nx��
_����	:�y�H��������r�Mt��v�tr��@]�������庚�����UZπc\�5�eMuO�g�8�����s%�,쩤*����4%�v�ϝ��[f��[()��߁H�;��"�ձN�7I��>�s�S���3bS�Tf�?��nՙ���E-L����6�����,e~�n`�	�çBxt�؄�6�Y�=����*7�� \΋����'��[>/�����e!W-j��`�ZM��
�n��%����Z�!yO"�Xx�����=��̒�g�N�hz��1XJ&�������V�ɍ�����[�T�P�dm���\��h|����"�f��?3B�14 �&g���@F)�Ӊ^�A��r���,�:X�Y�NnB<V��L�$�\��{z)(`�x���A�Ș�J�h:IA!�opi���=�wL� �
$��U� o`�L&Ub�H#4dT���I:_��Fc܅�'���zo�W���Я�*�֟��&DR�+�c�i�/��@e�?�K�($"ȣ�g����f&3C�+}��; �~�h]�P6�e�tD@v*੗�f;�bjV�N� ���"����~��F����d9a|nu,]7ʜ���rqcW�ɧ������r�7��k�q5BA9p���]'= ~�*�\�`k�T��F�"$��R���[�n+�F�d��O]��7Kܞ�2�=���2�ՠN9������aD��H]M�X��-���G��҉�|��4�oDL׍�NF��0�=u���p��o�r��5�����@0�(����U���Ɲ�B�f�����Z$�ݢo�N�]�^֩�;��]?[Q����,�=p@�@h��mEM)��Wj���������tU.q��0�LO�LV|=�Rd�+w�0���5W�?"A�ì�����xɿ���T]�W�AY�#�,��uݝ})���:*��xL��GA�i���֐�Ϟ1��Ŧ�"�3��6�� ��NҘ�j�a,3w2�z��q�K�:ـ�Wν@n�����W,�{�L�I���W�O���}�(F1�����tُ+�uB\�a�`[����s��F�mn���D7�`����^��ͧ�,�k�9�`�D���,Q�@�|�*��a�_�Uv8Da%�dv<8���{]�󠻛�U�F�Rޟ�}PB	��{R Iw�r�x��8��n;�@�Z�:�W���q���E$0-��.���V��:�����>fBc�$hM1����;�{
b�{��\m�V)�v(��6�j1��wEt��g�}�Mw�iR�.g>7#��XH�� ���i~0I��{�lm�8�:�ǥ�S|�a�u��~*8�N�c`�D�O��q+5S%	�"��T{k8i�n@'�t�9�iJ�z��%�H*�����s�<�h%��*]?()�RZ�/�J%�{��s��O)?*����x�w]���J^�d}���xG8�Ն(��Մ%�7��4rBSؼ#!��`&�0�3P5�N·�(h�e}.U[t�>Ў�r[[|�%�ۀQ��?c����`<�+�Ŏ���d���2�0�W9G�����R0 &7Ƅ�v-Vc��Sjt�ph�:���vo�VO�T�2i�~]H��Ov�My(��63ů`�;��&td�V�Y���4�_���2�2n�-^˂Z�M"�+��	�F���׫mCL��$���G�ױ�>'�4]:Ě�ja�\@5hu'��|E���"I��"�L+������@��ܳt���,�Lc�X�H�s��F?�T"�X�`�٘���=��2!y���_�^]H��c]��Z6����9�Y�k(����3ޱ�"���_5�}����*��4�E�4�^#
 .=9X�@�e;����x�۳E~�ۧ�,Kt:z[Pc��@��Q�X���c�sY NC���e:p��#O�8�j96��A��̭҉dȀ������N���h^-7����������֬9w� *i��#jP�s)А�l�qD�;:�1�p�N��� �UFȟa��q+3�a۷�բ����wO��O%���^�p�pu�/�(6��04���#������*�c�=a|�V&tuR)Vi0zbB��2
鄪$3�G�'�ɓpUN��4�뜏T���ۻ�=���<��Ns����8�&5���Sڕ�\An�qoN�&��KC۞7��B�Z8��]5=�d���%��4��j�|v� u���=	1J�v�H1�;��-���9�$�R�E���-w��\#?�4���'���[6�6DqK ��Z�r*a�ʹĸ�M�C�ج��R��u��yj�Ѧ�Ϙs������W�gG�~�J��I�K�VZ)<6���
�� [˂����h�����})n��	LfjXTuV�[�M�˞*=P��Av(��Ue{�e���s�3�s��f<�X�$�vw�����
��`8�S(pB���0!�(W�a�Y�)��Pw"��(��ޱ�������ӓts��R��)��=���[��%�C��Х��y��B��(jnqu�d֠����'J>��oV������6)_vS��t�����hӊ��$����~� ۏ�{;���ٽ����MT����Fhh��Y�3~
�*�Mn��Ru��*-�s�ITo�r�� ��~C���^��y���h}��k���j0�:��	{�V}�1R�ֿFCe��c�e�fj�g�$�;�1��mND�/�KoWK��	�[n�<Itz-F���]Jg��	R�&���	�#H�$�&�ar=���Js���\�d�H�S���
+q�l����R]�����r:�����b�}�q<�OSX�\�K��s���9���Dw�ʁr�c���^v�L:e�:[ZE�3_��')1��j�0|/�F�/t��Ғ^|ɋr��
fڠ97�vKaL'�����C�Q��P{䈯)0�?e��Ĵz3l���_+�	ݭ�݆��>M|TW6Xk����)������J�8�W�x蓸�g6�TD�SU9&�=2|��H�<&���5�����'W=�l�Gy�o�Qb1���ܳ,fR��P���rt�D��:�J�p�����8)d�J��'������ǜÕ1����{�Ճ`Q�=}��/���0y{�����%�Ud�%��$���kPUk���rB�R�lFU�O���}w�����G��#ܯ�Yi�`�z6�n�E��h�n�o�>m
�׵6H,����^]���P�f{�6�eJO��ec�ޮ�=v�{�r˃�Z��������hk@�s���R��W��mqVSP���>�"+ k��`	���Ja"�ͨ���c��f��x'�JU$�c^�[��>�2-TG�+�>�`O�E���>kp�g�x�H�V́�}؞�I�H�(���b(�8:�Z??l(���h�m�9��&H	��Q��\�������	:�c��x?��S@Y��㶠>D(�AS�o�+�6��s-m �==BIWZ��ź�W�Hxۏ��ۮ!�e�X��#�)���Ӹ����ד2+O��v�x;���DxeJ���V���G���eO�֚�{�s�SH|;Q�MY����؉���!�`������y�X��1�o�4}�4a�K]��i���z瓤e��ߕ�d��]4C
2oʶŐ��2���s�t��m�yI�����Ӟ����)�
 ˻?���"l�@�"�h��|��E�xB���E�ԕқA�k�sk��x0<V�a�)
�l[VP���r���Z
�޵�3�iq,�+?��}���P��?VOXb�y���`��Yp�:3mk7���w�'��C H��g�=F"D���`0�v���!h�����q�)UE���B3���G|�~��8��� ��E�O�,L�I7��N�� ���Pm�>�z
eH�8����Lo� ��p4_4���c]�L�z��&���5�0�Fn��������rQ��s��W.�b������ͫꯗ����#`p�t7�q`Q%�u✅�V��oY�"����Rb�4Scx�H^��>]��s� �Ȝ�\�x�Z����OV�;�e��]���3�orp(��҇�� ��R�Cq��:� ����n?��#�:�גz�*�̑@���go��� !��r�=SbK�n`��^ 5Q��.���o�ܷ,e^�0��Ɩ-$d�?��c!TL�	����Gj���.:��X�����?~�;ջ�?������V�8%e��7�^���������(�Ԭx3���g�=��(�_6�ڨ7�	���Kq��Y���,�Rv��MN��U�f�Z�;x��r�ad=���a���`�6�M{��uȿ�Ǥ��n&�ک�:ڻ-��O/o����td���l�\�Qk{5)La�ـu�ف���u��i��)�Z"�-WX��c�$5�+d
�:U)���L-���@}��EK���0,���zA��Pǎ:�˱�s�\~ď�D),�E�_���n��C#���F�_,�0���&�Aõ�puC�^��J�]"�,�`lc�\����L���k�쉤���)�&�c��������L
�5�
گ�ȚJ�F\�1	�!�5YJ���y(�S:��f�Rc�\#R���h��8�eގ�p��M�ޏ?��O�3�Y���0�!�x����A�U>wQ̘��7�r�cmB#�ʩ� �]��`�N���? �R�Zf�E�5n�$�O�W)Vי����H/�Eh)D�k��"/�����^�E-�XU�.l��ws1Ⱥc��]�y�6�%Ft��x�&~=�Ƿ'�Vs6����]���uU?X��c���Eb����몆WY����~��,�{g@��%3Ɨ�����ַxm���������p`�XͤUE����5f�d�(=��kdmn�+S�'15��N���w��������ezqrا�z֏؜�	�o�O�{5�Ѫ���ЖI��aʎN���nXE�8�E�:��+֗�C�� o+3}�>�S�!����W^;�Vy��d��~/>؎T���'\�nFL� !y��C�Mjof]����2�c<�����/m�3�f���a�B�5�;�ki�Ij��c���.�>�
7�R�}�\58B3[�t�f�ڏ!��">5��u��,�����i5Z��~F����V���<	���	��w��t1O�������̮�e�'w-�x^��_F�7�����ѓc�/u>��a,{�}{�c�k<c���CM�M��+�����j]�n�g���+\o���������f���!Bc���S]ʯ�@bE��?$�	�i%(��Os:��(��p���-[u�av����$���s����eC��b9���I�L*�&�!����+� |-~�,1:T�����O5Sg�Gd�oj�n�MR܀�ۢ�i�~�~Zj{h1�X�bN*<c��I��@�ޡ�H�	��<�b��(���3�{₲B��[�n���峘r��H�����.�4ݓ)G+��_A1�!w�7�Q�-��o����%�K����:��*n£:�6"���&r��ٌ��  �þJ2�i���Q�2��;.�eN�
�$���=7��F�H#�L�,"��D$�yW��j�(gv�ז�>R`����6���Ԏ�����u+�=��x�F\�By�e�H�%�q���1F�v�}c�����h����؇�rgz��9�����6�!EX%�~J���ô��Bs�[���.c�n$�6ڳY�Ƙ��m"V��-a&��������;�D�H��L|�c{]C��([ˍ�T��$���c�s��y�^��F�C߅cLa	/� �?#dU��pn(����J�k�Xd��b��ޤ�@���no+���+�_�dI�r_�L5�_D���
���z�ɏH͓OHK���\�C�{�`������n��<�; V"�N���v
�"Z�ݮ�����P���E?������$�6l�S��/,�� z4ղq`]��1�L7�V<CS"�8�k���s��J��:hvu�c'\8���՛�����Ա��f
�uu?z-�2\ɇz)�m>'���tH7�RA��MW|Y&߻�H���$�X,�
KL�Xk7�2�f�!C#����C�x��Dӻ�F����˅3aI�R��)�����KV�H4����\{��5\R�g�����wV0Q�4�`���)x��c ������,|�7��3�]�1����N�T A�'�HZxW�x��Aʨ?N,&5K2iE���P�#^J��9�� ����.%��QLIP�k�TC혴�gTɊ-���WɄL�!P�h�ç�C2]k)��]_Zr��u�5���]��l���G:��w\�wh�W�K8��
��>7A�s�G̐��^��^��޿�)�>]�,N��7C��Z���Xz�f#�9n�����"�.��K��xg�%�y�r����ſ��⨾��'˼x�'<ҋ��B���/�Oᄶ��S�?t��Sr;�Bp�E��-����N+Q�����c����>R�!�m�"1��l�.v�57.�"��t@�D~a��-à�0�[��,�*�࣠��jH���Q] �.p�m,e���)Xh��)�/�����KI�W��u#���L��k4&'�g��&S�V(@a+7��j��.��k?��L��鵜��@5$�4��1p�K���-�j96�gK�)��I��m'���6��T#:�_�&�W%�A�G0n�Q��q�����.��_��ϏE7��*���Dj:)����s�aJu��P��u,I��Q�)��z�<�b����j>��&ξ5�VIөwI�AdA]��y�.Ӆ��֍̋����#�OUfw6�,N�nt�O@��\g�-'#��[ą2��l�5�ӔZ��ɏWT�����ۦ��	��!V��j���B{]�|6��-����c�d��R�j4;��ҹFEPQ�vŊ����7m"1R���B�yO�n�$�i��:ՐmO H����������i_�u>V���b5.ti�{H�T*s��݀�!#�%�Ⱦ��Qو\�SE1���]��	��y�NB��6r뇫�L��sӬ*� �u3�e��3�O��
Y,�>��W�7�89X�H�Dd�'�ʆ����Մnjp.�;��9~���$��}�"TDP�i����!���	�{hK�_J(f��mU-�6����q��*���%�cjq����G�6ӒK�;iZ�2*�L�Gw
�p��`m���a�BQ]QJ��>��1R�����5`�N5\�;$T��k'�7d��`�RG��l)1�'�Wm�%��x�귵����k��ô\Q^EV�KƂ-�����H��4�[�T�o����k�M6�Ρ�)�gjΕ�T��e�o'�8���|\����dC���l�xdp��S�4䛡o1!�����\��M�9I����q�	� �mN�J�50/r$g���h�DS���5 f@���3잍W�w�h*�8`T�BM�$߱]B�@��W��ge������Lg�O�'}ǄF���;�
����j�k6�[E�����wK�c�ʜ.��"kK;B+�(HiJՠQG��@�rj�����)(vs����wg1���m�f�Vy�	�d��*��o���M��1�w�񉫠��Ҋ�˞+��9
��TZ��bsb�*�mt|'��	A��6�N��q���և��S�&9I9���O��`F[��?��W�����NCWA�IC�6��b�9?��,(�d�w����
&gVz	H9�V�Mƅ��z�^����
r�DI�i��ީ
�u�m�)� ����?�V`R-�)����0TS�1� @�Q��S����ڈŇ�k��;���/{T��L��&EX��-�,l�/DK���3{��E���>;(f'��oJ��	���}�bwki�.M�~3a�;������x��]|2�wT�T�"���=���hu���xˡx=i-Mt�h�0����{Yw����u,������fscI&���B$}���=��U�m�&»���XK�����_�k�{����w��2W�s��`�6+��xA��i�'����as��FÂ����iܛ���*�N��,�%1����PjBr'na�W�}.�٣��z8�3�aFVXG__�,w1��>��dKu��	-��,>�9<����A��J�}�!x�+�T��@�W7���Ą��-���Ƭ@�(��]d*U��&� �V>q7T���Wc�I�xh(��g�Lp����Pq��r��Fg�^ˡXD[�W�c�#	΍�V"[�͸:�0q�P�[�!:pŝ��6���i�U���"��!_�j�����H{�g������8q���W�0�1�m���V�Pkp#�C���U4��U&�^�l�|�J7�����:G���R��CRR�,5�t�����W]b�$�,&}ϰ��y�WC�qc>
��e���  �L�"Ju��o��l]cn{.�e�$�X).]�Gj5AQ���l��h�{ő�wc	�dK%�rJ}K(�b؞�9��v��6�P1���]B�=̺\0��~���/�Qۿ��w0�Hک�܇,8�d�L�X#x�|���1�7�����ǣ����y���dd�^ԐR��F���o������2[�S��O,�UhZ������+~�9��Z���9��dI#^j	λoTΎW��*���Y; �ж�Jˤ0d�U	4BX Ƞ�"܂0=� Y�Qک�n��L����b��;5>4���浮H2�N`-f�s(0��HIޯ_���v/�#C�H��,L��ԑj*E��q��"�IR%w�^����Ĉ���CKyq^�c&L70�^� !�<��5d�D�b��M7�ycZ[?C% z����+/�#?1�GQ��e�cR��W�o�;ٶ�zX���M����A�����9��S����w
�b�_]K�y�ks���bm."]���;�|�Rޤ!�S��[5.r����aZK�H��@F���\�F��)oZ���k
�U���9k,�zLX��T��j����?���ƀ&}���%�/��<ʔq��٥�o�� /`4H�㽱튚��
֦iUإNl�lfu�>ص#�LȾ5�:��в�7ꃐO�����H�vȨ:�����6c_�v�{�ױ:���]z��sɊ�_��)�s�����sIfZ�,�5ɵ,��g�	��m�J��7b���h�/M7��M�a�zQ,`��T��!;�eJ7�)�@���D5z6�Q��n�?�!����/eFrc���X�K�q"���n`��&P��F�6�c�Dbl*:�c�e��ъ�HwD�4���(��:gd8��{e��j�=�pݣv��䊱+nB"L��[t~�@L����˜��z��f�!ȁ�b�E�㶩:�M�޺�>��ﮄr�<�E�MEL�}}청���
ه_�*d���WB�]B�$s�p�+|�?Қw*�)Q�>E��6yW9#BSX���.�H�����]��7�h�n!���J��P�O�D�:���T6v��D�{�jy���&�m�YeY�_o���IzH��*h�?�xI���V����_0�W����u�5&ڍ{yF.Ǡ���g'�>9�-4� �ai�ɷ >���}�²
_��O �����0T�<+LW����	����g bB�'e×���}���hq'���#�Z�����@�E3���s�����q�����<mj�6�B�є;�[��́a��db���w��}1�����J�p`��M*�)a�]������sӛzXң�JM�x�@%b\N��%#���{KV�::�t4��G���I0v���%c� �9o{���bM���nyoLA|�x�K�4�SH���i���]�ܔΔ�91aQ�A.��D���3n1�:`)�X�k�x�@4�x�W�8�6� �ǒ�`U˒��	�F�X+���3�d�I�#1	b��i����)�����.��Fm#.wKI03��o��%�W5��8aBv�š/�C��mtT�o�vSQf�h>�2Y���:쌣�ETGc&�͵��p�P5\���j�cr �/X�(�" �����D:���lX*Qո�5�{;�"�7jȿ�&��4����S�Uѻ�@o'�*+�:H���w���`�#=����H�ބ��˄�x~&���Tco�/�����t�^-�js֦���h�#c�����#+dx�q�6Z��X��Q���V9��l�6��K��O�n�:���˟$52'Ꙍ�ۜb��C{Aq����Ɠ��W�x��E���GP�g��+ߺ	���1��Y'��3�}f&A���B�vˣ�.�D&O�M�RZ�W����1�@F��*�'����Γ=�~å�3ͫ�"�"��`���o{M0B��o��.m@V��E^��P�gm�}?~��'�Z� ^�k	�=�o4#�[�x���/F�	p"D�'�c�qD�u�"W��=��A8��IEی��4�4]kQ��$�1#�v}D�]�FYq��B��x]x;�./<2 7A��à�HP�D �k�+�W�*���k�t>�(��žɾ{���+�5�xB@F'�Z�g�PQɻ��|���,2�c@���Q1h���7�-��+s��?>b�քoy�9�I:��rB��� 
��O�.��wh�)���?��"e�}� H�s��9}����Ô��2N�1ՉD{�"ϥB�. � _;$�D��!8�u�^���l������|�I�Ώ\�G��u���Mh(ܦ���+rSV擝
���}���|K��@v"�ǌ:3��n�u�[�zƴ�>�;�4�9ey�_����@��_���b�wa}���)MAҜ���sbٞ��a	��9��-Ŧ���5䣶"!d(p7O��[�����ތ���4�|�7��t]ǹ��[*k?��.�V�2�`J�}� ��s[��O<��1�wy�&�0�J뒱Z��$9&���8t��v��#S��LQ��4�b�� v	YS�/DJ%�d� �o�r�m/�b�F��u���V�Eq���T�"%G#?x��|����J��"6�U�,���pg���,���9nx�t�CO<�gn`P�S�Y���,�5;�������ۛ�&i��a��>`s�i��l�PV�O�M��ڰ�a�t�(��^�8*�Rl~���B��"1�6��+e�TOϦ�D�����Ѝ(A�����<(,�/}��:��qR4k��j��)GH�������n��$~G�u����\37�U��Y�M�R#O̦�� �[��B���[���j3=_q-��9��vk�y�S,i���Ǭ���W7�jh��	c��!a�۳9��U��>S���W]v/t �=S+U�3m^(�4��lɑ�7�ft�]d��)��xPU��d�	H����T��<::�(����jq�]�����a5l�ٷ7��SF�҃P���"`Nu<OF�����=\�踐�C�-Xa9T'68�mJ�m^��x��̀k�̝�� 8������b�/������;J"${�lV�&�����E��Q{�=m�y-���? 6%�`�i_m&��+fA&�Ѯ�mMwdG�Y	0�p�[X�ܐH�]��UE��*3�͍W{�<5�]iw6��R���9���`�*їA�O;�O�~#�s�a.|`s���
���8vg��#�eF$�⹍����˲��� ��[��HV��Dk	��,���/��3�b�M����U��yV0oW�&�eDd�q�!@�[uv\u�ں��U���Dj�F��:P9}�N���T�s'
g�������2�%���G���J�"a�����=�fm������H�/[�Y��áo@�)���F�P;(���kע�Ms�0��e�<�{�2����D�3�iR4`l��3�4���3�i^>AR���z��2�V�"�E��_}�NlÙ"�}��M��x0� ��P�q��!~��unҺ�aP#@���=��E<uu��E�X"7�q��j�<j6PF��3��?������t����=Dw�	Q(��0�邥�g�,�Ů=t*	:�
�.�>��a��1S?�s�Gd��Y�β���R��|��O3قB�/�����T
�#'՞T���X��I��&�>����+6�v�},v��u-rFxz<��N�!R���S~s+����[�	�M�OK�&f=<ζh�ʕ�O*���=r����h�ħ&X��쿄*�eږK�M��̗Sc��'!au�kͷ�KR��^^��GK��~t�W�����R?v����ޅ:>-�;ύD�
Ɇ=������6�!��ǈe��'��آP��A6��fV�ȋ8x70l>�$��I��|�	u �A�F^�(ˏѼ�ߖ��g嶑�9��s̰�xx�:����Z�I|*bbq��⚾�Zz"
y�`����;�9�&yS~a�ќ��X-��?䘳���͹��*��� ��ğ�� �Ha� &d��	��0"u����w�Q��@���Lg/�����
<o���D2��Z(�{Q�4�I�l��|�bD>���y.�ʍ_+�\�o�$��.�|\�𿺚S�4Ǧo������i�$>]ZRn��l-q�J���&��AH:5�/-�o���K���������O�MM�l�l��HA�94�;�zĵ���P�$����n�Q
�������۴�`XU�+{�/�I���+5]����+LO4}A�i,d��9���'h�R��l�����og��6*�J�s�$}���a^a�{[{SQ���1�1��9�O�UuX%lf��t43������h�/�wq�ؾn+kP�f%�V���dK�6�a�Tʢ5�f�qJ�L�^df��f#lz�{�M��Å�r��=�*��6%��,��-E�B�~�i�\C�P��r��� ��n-��h��_ԃAav��v�E��h����J�hP»���1�������"�K(3��Bކެs6�֕}�&G�τPw6�y��\�nX�w�Os���o�%��q%���Q�6����!���k��V�z������- ވ!�*���TCQ������=�)��,�K���R	a�Ԥ��Ӱ���h��5�U��/O.�>T��7@�gETߺ��ٰt�ѓ�	�6F� "U�O�/s����aһ��������kx����ƴO~��I�Ó�����]��~7��e-j/,X$��c�:�=��tֺ�j^���+�o2+v�3,�縕�����J���i��R��p����<g�^9Yl|;���0����ا�_01�?�� +���U�7���h�Q�h�I��(Z |6���O��C��?�:�cˡ��ei7~�&)��҇�ns�Q����6��K�1�+|~�^��+@ph`ኑ��3זu����K�En��e�Ƹ� AJs0��W���
�N���9�uF�N(�[��w~������Pk�_�O؅�Uy��u�����x��\mJ��xs���hݒ�蠳�&'X�__
;[���&�A��r�!�5�c��@�Tm���э�3������H. X���"�n
��	�����Ij�2�>����}pH�S�(6����=��?&	7�W�>ROf�D��L>�w(>h\�R�=WSoSO��S'J�_Y��JL��V,i$��&i`��[bER?f���谼?��|��U��+a�K)q�r���Q�Pᇲ��~��n���S��K���q�[_Hh��]M�D�W�?q��~����B݌�w��À�P}�y�<���X���J+�n���^��h�5�U��ϱ����:�1����A�Fɕ���A�2e�o�^d�](����nB��3Е�4����� ���3ح9����惡uQ��%��P�޽9�Р.�tT�EL�I���Kǆ}�[�O��ɺ3B�v�x�7�VZR`T����U�m8�a8���$��!�o��6a�c`$	�+�T
 ;>��JV�K�
vlפ`�	�Lq��_-�{�BM�(y[rF�(:�ϑ�3�#���|�ƀh���0�����v艩9�~�zpU�5�.�Te�@
M�1;��WF��iOYs� c]���� 6���5g���Ϛ��,u�� �t����xe����暴xl�i�Yj	�[-�V�f&�s3�jx�<�0��mpǕ0�m�_�]O>ڝ�m��M��G�W��2S ��h��#	�0Ƌ��ћ���o*B2ĺ�8B�F�d�/�,58Cq��k��u��w�'�A����7�v��e��ҽ�|UD	׭�lZFD��fq39�s"�{�=[��#�R���L��&��-G6]��O'�iI�O<��ޣE�i����ѲV�l�H�����?F�.�c�.[�d�-� B'C��Je��N��قx(�
�1R�q�WC����W��C����[t}��
16E�w$`B�<�[����
�����d��a�PAg��$|�֨��(������o
4j�H"H��P	'b����̑�%�V?�K��}Wέ�Н�9�4�Q�&��t�z���ew�`�΄ �yN,��[mY�l �V
!}^/��[E��q�M@��<�|k
%:Ӡ?��/�� �x�iR �bm�Fd/�)�H�uY�0�?�׾�(���,J׵���|�f��d��]j����$�OD٠��73�즴�C����/�Y8���2�d��B$A�UUd2�
