��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU����ax���Q����.�Ā��{��𿅍�C�R}pz�^Kl38���]�^�V!
�+�Z�	%��M��L�~�����9G�*)#��t�c>��k�rpP$�W9[����jK�����,������7R���>b9���c9x�)=���-qS��M�^Y�� �ޒa��	���'�Y04�DW�[33s�PWXn��7��"��u��s�8~�0����y�d�#�`����_�K�Ա/ �ݍ<�Sq���J��F����yT�W�r(C"� ��1'0� ��u��d	�Ԁ�y����$���Ⱦ�fE`��B��O��4�4e@݉y�O^����t�_�,�Q0Z.ۯ� ��Ii𨀱���n�eSy�AO=$�9�Q`���5��P^x�������S��[&����]�2�2���|��bS�.ɡ_�<�X�-��ɀ*|9��(����A������4��1I�ϤX���^�����JR�Y��NA��.��WAn�DIw���k�֙<�|pC�h����MHk60A����Ij�BB���\�nǾR���������r,���^��e g�6\=�	�jV���sEQ�і;�1M�a�Ld5��AK��ͧ[��p�6�/��z:b��vÚ�pz&Q����tf�C,I�W���H"�|�����`�[u#O�k���h��T{���5�x>�K	���O�����8d�N5�w�(K�����C���YpuD#�V��6���^*�B���t��0�����\9!��Q m�wMQ�Ml���zʧ�k�Y��|>bF�-��Y�ūM8rC��o~�a�����r�?������ M1!�&�A�,/��
15��4��z���j��Pw���b��|�Ӫ]+:1�q�/Pmb��C�dP�)R��6ɕ�&�%뿀bɪ����q�x_ ,�ٶ�*�!q����Xd�~�Am�@50l
A1D���g��_�:��on������ �8�R�I��s�b]��IP��4��� _f��_�n�}�ӕ�W��ܩ�3K36�y5-=�E񹋰t.�MR�����"���<)�>hj'����Q9��^�g��O.H*ˤ���"�T���-`�m�[]r�U��;�>@)bUC�1*�U[D>�w�#�Ҝk�>�٠ ���g/w�+�&���CYޏ~q͉W�to�?I�m%�B����ܷ�֔��Z|{���n	����$�9> 'D�ҷyo���k����la���,3�OC��+U�E��Ӗ%��>���%�0��?��ք��}:b� Ɗ��3�;�E�IC����|�+�΄`R�:�T&�6�2@��.�,Pi�0	�l5:�9���g��U���hQ	X�����yo���(�Vl�Ꞷ4���?d�0�)���)/4��ǵ��s��2�PQ��m�(p��� e޿�1Ŀ���,"<�F���3��H����*����oiv�8T���)
�9�_X�l|s�6�Tĵ���F{�}�:��Ҭ�d��m��7��!ΏZ��G�ֈ%��/N�Ϫr~�,����<+����-��};�Z�^�	�٩���q;�;�D�y�B�jd�����]+�� #�`���{��*P�p��öK��!�w��`��t�i��`�O���	���jp^��3aZ��T��[�`N������0韡�R�G�isR���5H���c�3 CB��8k]�aLNm}�(e�l�B�z0�;+��ҿ�Og6�t�f+��U��;�K`�����M=�I����C������L�h���܉{6�L��S�eζ�8�u�3 ���-F=r��I�މ��R�_�
��?(�e��f�ط��.u����1fo�����Z5�Pa�В zɗ*�|�T�Wd�D�_+憢�Lv)�8�q��#�k=zQU��P���p菊GAlR�6<Q�v�{�,�D�:A����1F�!7 ���}4|�%d����loYu�l)��sZ<
`��c��������+��\[�&zx�i2�#�0���E����c��okz�_�e =Շ4��p�J�S�2���Ά�$5q��¶+���	�0ߑ��؎dpe�-�h���tr)J(��+&���<E�)!���(�qy��6/��R����g��C6] �k�B�i�)�pB���'��vJ޼e�T #L���M��5�m��&|t	�A�"(O�H�IF~B�*}�܃]C����QsA���B���vF�m�<y�q��L6k$#�d&,޽��=�1U�\�f�Y�y{2�w�� Rz`H<�ڴ����뙂z���ZXN��rXW���j��T���'��렟����\5�rxkx�q�iΞ�)ŷR6ʵ��/�%��<��Ob�L}@y���QD�M�%�ǔ	��HP@���Xth��k �1�c�G`i%�rl�B)rg�{�)�^�N�?�Ј�WR�"Pt�i�'��I���$��%qǛYƉ<��V༼K�����A�l��XV�v�gI���<���ٚ�����)�޻�\���A��5�&xe��q#�ZTc�Yd��3Ŋ^eA��Gy�4v*���6]ߨ�8�tU��v?�Hr$������J�iR�#�o�b1���%�X���&��$�Q�;6���ƶ}�#8��O�m�䘾��q�_�W����҆������}D��K^�I���/�:��-*!�N��S���靚�Ld�w :�(g2~D�J�Պ�+�2M�P�Db?��x�>\FxW4z�M�f�&��m��`,��|r� �n��	g �y��x����;����{�շ[��L������op%|�����`EW�������xwS)�����z!	�fl��@_�1'���3�����H���^�o���Y:�Y�X1�-�
�on����[v0Y��vo�~�337�g�<�ʘ���}�b2�B�#A0%fP\8���������|��J�U$EŹbT�H;�R��_3)��G����w��8jm;�3->�[Ā6�c l�i����Y��fț�۞��zS�U� f��Oq�P9#����b?H�J7��9���&�S}�u�)�F�Yk���A�� ��t:cJ�$F0��by����멤`�,��]�V�*�<�A�R
�Ϭq.7��s�J[�RRWi�	�T���E��}J�fyü��Ln���Q�� [�/eP�%c�&�m�	'�6L���sxgs��ӛ�Y|���tYoS"�bGD��h�d��}*u��I!���e��	"J��)�>��<LM]o����l���][kf o�黊֡6R2�~G`v�h�d)Ξ��TR�����n	7aD��V��K�!H������o��w�:��՘�6�Q3 �X��F�	0,�n�p�x�lh�SKF��%������62��s:���D��`tQ�!�.�za��x�+�?��-!��.��� r�`A{�n�=nV��7;i�A3����K�pB�Sm��ꎀ��u�T%��2�V:��L
����$5���dEA�Ɇ�˙�cG�6%?�(�W����u"��˴;i�����m�J/)�BH͡��a|kT�(S!��}3W����Y,��5_�'�6��ZSk�xN��"���즎�\v���������
uSf;�~,H)g���FF�h�L�M��h�!|sP�?���[Ն���E��X?�+�?��V�N�����R�������I\����l4�:�BkJ�*(�N�5��-��a�q�|�Q�Ut�jR�:�����>=�
#>~]ac-^[�(�*�����vg��ԩ��3#I*akF�U*?�֩�Ѭ�����z�-���`����
�EB�b<���t��+y��wn�b���T?��6���$�:����b�����NliR~����f�S��qσʘm7q�+$�``*��,%���}�7��5A��c�z�Mg~ij���.��>�N�Z��^�d�~K��/�2��HQ�q�OU_`5��vVۧ"�Kw`��vb_f��<�(Y����R*Q�#��� @�x���'���Sb7І9s���\�}ђͭ����ҹ(�T���U�B��w��,�Ds/ud�$N&,n��q���d{������1����ɴ�IQ-��+�u�8^oK��1�Q>4�-���DBE6J�}�P����+1����:&©���6�<ϥUu����@C�r8L�k��[�7|�0a�:GO%�Ǉݚ�u��?��j��4>ݶ��}g���ߴC�Eʷ�(׳	񇫎.�Lo�*�֓�E�$+�5wE\��Y?�죶��МE�?П�F��|�@�o���O�3������~�GN�d��X>U-��Vv�������;��%*��?D�,�3-���{c�a����ѓc@�*�����ll䵞W�yt�%H���d�jݲ���O���^�s�q~fԃ0�<gE���$���e�6�A��m���Q���t�9�}7�����7��a���Jq��~���6�㻈�5��/?1o�����'W�SF���@�;����zҒ�O��J�������>����W �al�W���E���\��s�:p�v�����5�#m�t�t��JL����Kv6<|��r��P,������?�2�Q�rkb�4�bVn[�o��;��>$[)��/-�(�):�������wiX�N�����$�G��L�hZ�1��2�3aUv�d����\Y'1� �\͌��+�׈u8H/>ܜn��d�l|F�u	tnKx�1�7�F������JP6/�*̧�o1�YEa��p�� �ū�KTPU�Yu��-��Mr�.��R#��j��o�4�h����2��?�AA;_7�Jd{�`i3RD��SA�X��^��K?���#{ǭ�[gtzˤt�]�D��B�D�jF���3C	��)�K���S�ł6G�6"�C)��2<�]����0��V��nxbM�q��5�E���a�L�$ehd�EC�_9��<xUp���/�&�a}��	�Bʗ"9�u���[0\�ce�?�2�h�����ӡ�##��A?F����p�k�ly<�a���G��4A�3�/�c�#)��υ����F����׫`��-��ȼ0V�uM0�h�-������T�gy��qE�b��B<��_��P�Gaڽ�E�����q�u�*��_�#kU�1դ��4%ؠbI�2��f:���KN���윏	�����اfճP�� ����3� �����\f��PTJ;~���9���Y)��>��$7�i�u-�u��mQ���RU>r#�L:}l��bbl�����d'�B��0�؝>"i����i�������d�nT �P^�{8����)��o,B*���G���E^����>N��>�}e�LX�H[�;�UUiZN��~ĕ�4퐌E����u�Y���S���{��c�D໌���^�6k��~g��gx�H�*���]F,A��֫
�hx�vb�&q��`��`����ِ{*���f�������Ⳉ%���2Q�<�̪���yi U��T��'�� ",�)��/0}&��#� ��
�	�X����qm7��q驥d�?In�RN!#���A�|�]���E���4��a�c�>���87$��m:QﴣQ�O�։��/��SQ��5	����jT�"��6�^MD;�gG�|���]��'_���H�D�����"���cO��ڠ�"���DΡ�]c>�n�9];�xAE�6õY�p���2��lr㩕��R��U��T�l�ڌ����6(���+���~��s�N��o�o�l�����~ފR[{Da��˭i��3���ߴ�i�Q�7 ��9�6ᾓU���7e����k�j=�
��������ccp�Z�"��C�! U����Mۆq�y7�lUIP�-
�C�p�G�ý@�̤��b�XG�L8OO.{lֵ) �[\�⼭��>�p�٤���5�3�Y�7�P��C��v�R5ΧD�
���ｎ���t�!�һ�<f¿�a��55����&>A�ef�]4a��˛��!S��J�!�hMɂ|��^Jqv���������� j��RW��A��a:6��'p	0���r����Qyx�i",)����^篓����;p0wy��ϲ�ڭ� *����֎F\`[�K�qʴU��Y��"+d8�f�@����_7�@P���@Z>O�A­�_�p8L��?�< �7<�`������A�ܲ��k00$�����p+@6���L�ʪI4���d���$�$7Gq��pw���lG4h�p��/����Sa�{(�z�J�������8e��pZ�C)��"���s�ӭ��!I����ֵ�͑}u�u+�t�cs�M�y۱�$ �s�A��tqD�t��hD�s |�4��Q�&�Ia�q
ېT\k��[�U�HOհ�����OJV&�<3����h�������B��$t��vb���A�9��.�ơtQ]�٣+��%(���=��z�d��R V�F�%��@8����.T&����O�+K�)L�"]��|�,e9���O|̱li��@�/�����Hu�h�{��b�Dcs6��鯼�>=V�Z��]��g6���xV�/c�ʑ'��Bܾ��כ�0�G���[L���6o*�v�oor���c�%�oII*9{�j�ݯ���no�[������]	,�9��hO�Eҗ����j�����'��&���������cӛ�Y���B�����d� �	m��H�<4V�Xo£���Ѕlf'|�Dl��k>X�_����̙p["�\&�1=��Crw;|���_U���(���
�v��w{;8��	sX��^�/R�LԦW�Dn�}��3u�o!�\d��(�_���x7N�B]Wu�����͝�^�X�����Vw� ���ܓV9�S$���<���m�����E�l��yR���ƚgk�����܋�c>��4��E�]n��]��H��!/�B��k ����d�
&�ƪ���.�nf(���§+�9�9~��q���(^�e��A��y��+�T;��}��S�>��(�6ݷ�_�ƃo���$@��1�*˃Vu��*��F��E��+��MؽW�Y^�3�`,y�'���-<��?fW�+ ��%����83v��.������]u6a	<"��x�	D��qO�Ι�@V����F_��N��`7����j=t#�,�ڲ�$��� ʑ\F×[~d>��D_;ʊ��40�T-y'ĵ�ы���	�fZ|M��^��G3�3��3��1�+�֠��	��;^��M_(Y��&'�p����B�����[�ן�<�*�� �c�_(�k-��!s�,?��FHT�K��]���:lK?���@��MV�~��t.�(���n�v�'f�Ni֝�`9n6���{z����@��w�5��,w@$kk�k��}��e�)���e�86"�`b�vŇ��U1(�~F�i�E��x�1�<���5�E-l��I���m5g!�������Ͳm�:�P֌h\dԼ�ڶ��D���ǽ��A�)����` ]��Wf�V7&�FقΟ�K�٢)�LO�*(��G�PH�0TY�4��mߒԫ����#v��|m�{�U��z]qdp�0LX� ��뀫���/ vi��L�?:C���A�"�?��#?���*�7����J8��J�N��.�rs4�q�;�I�$����T)O�7��r�M�jyb�\2K|�S?�X8F���m6x�� ���/�i�3�`C�Z�KG[`�ӯ�/�F=˼�z>�ho��M��b^��e�͆iC�5�ɏ�wuVh�C�V'�Q��=��^o�m$v����y�|�u&)Yw�L�5S�Y[�����/z��jf�O�N�f�TZ�:T��t���mfn�+&�s��Tn}�D�����Q��g,��oI�J�-?c���hʒ�Y���/:49˃��3}��m`bܼʓ
��>�8���$��'o�b��E�۷�b��/f�8J�> �����,������ˈ&���C�[�����Bg��Z�Y0���U@�X,�i2���·��!�� ���f�R��U��C���fi��x�\AS
�W��1��=�����l�a�L�;��7�t�@��D�/ȃ���oL4MX�����@&.0����4�QzE'��_�M�[obY���h�t�Ԭ����)���S:�R��TP���FnŲu+�1�P�3�vQ(&�X��vx+f�2PJ���,-��f�d�����H�"�/�'`��̫��	W!x�x9i�a���KI���E&@" �j�7oR�$`�q;sD*�K�g6 C�@RI���F��Wܴ �uH8䔈��l��6d�6H��5QcȊ��3RGu�����+=�3]���K�<��h��D7�oϱ��pg�{	q�GnM��yۨ&��pq��\x���6V��vG���ԕ�`����N��a5�������{������t�E8#�ߒ���%ޏ�7��� d�Cmt��@L�+�#�Zm(Ԑ�ss�)�����#�������ujt���w���+a�LT��(Cg�} �@��K���ʵߍ�>)r��z��f���w1��`4y���Z�H��Xxox&�.�!
(��7��g�Q����xNv3�¼��P�9䣴���{̇�;�.�U�0��<�iw�写][�>VA�$�QY��<~�*���6;+	��w̵H5�$d�s�v����}Z"n�t�|�4Z,� ��)��N�wQK�r��P�3M���3h�뽷ĕ�/��--$�� ����Ф��Lj{>��"lU�����`�q����Z�+1�d1�BT�ؓ���{PX�q�M�.x͖�Cjr���	��v�&\���雓0Sx�%�n?���b.�BX�E�{��Se{C��f�3eƈ{ׂI�/���lϩ����l��]7����µ9�W"2UG�Vv����f�bP}�Q����E�����z���+�d��X5f�_1]��jj��a�[
��"����Ko�)B;� .�@��{Z%v*s�����%P��A��mY6��\�/7}b�͔t�\��,�^�D�x�E03��ޒc�L�r���+�:ܑC�%��$ծ(L�\Q Qj@�t�-[���\B���A�*J�4J����Y�ҩ?��5���/�!o 0)2���'�����#���x|������%S�a�d@�쉣�F��������>�8F��"j:Y���N��Q�1K�i�9�dڜ�6��_�x������u9�㇛d�!*�Sd�&��C��8��o���\R9'� Э�$^:dҨ�h԰���9v�=Y P~�A��Bcr;������'�������ea*v }d��K���;������۹�8}ea�5]�>���T���i��u�ό�h+�db�	�\��}� �}����Ζ�\hK��/����;\]x�$5�#M�S*x��<T�,U����m^x�CN���x���� Me<��[�@�?:�V]Z�KH����o�"�/�Q�;��ײI�b4T�v�x^ ��`��
�b���zm+�,�A�B1(�ȃ\]J��>��D��Y-d��$%�f��#�)���g#f\�z�x���|=M,�2�W�d��� ��D����l�.�����!��'� 5/�����3����W��4]҄�{��g��ˆ�����y�����E�" f|��
�+��6��5qJ�; ��|�| (G�۬O��Z�M�� ��ǼW�|��Gz�2o�q��:����<��,�-c�,������8�>�u��)٨d��?tU翬�&e��I����t���.R�;�d0yl��-��	���JO�'b��f�Z��u����d�@��W�"CX�X.���;�&eQ�/׎����v����2�*ݦ$�GME&�dV�.ˬ:�����AQӄ5ً��3�����y�]/��ܻ8RF�|�!t�kiO��M�|m�do\p��ɏ��<���k�H� ɪ�v����pp�,�n�J&���0t$���v�����MP�1�(`T`>pB�����|��E(��[n9��^�;�%z
~'�e�
