��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��2g{p2]H1.3��{0����E��&I�}ԫ>�2ߝ*�1��\u��W$8�M�"jckpI	bg�ËF�t�Qӽ���%�����Z)�S[,Ưe�"KPـ��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��9V�H�YpF�t ����6�hhu�81`^k��'N�ȉ�p�A�V��/�^�dl,V�_�$(g���ð,2��i�-0������1`!y���X�!��!���p-���������$O���\�P!~l�̡Z�,��l޽�E)���R���Y�q�'��@)4<G�X�IJ��e1;	J���?6�{z��g-ʗ)��
E���
Wk��G>�dSi]dSɬ���9���*d��8�[{@ھ��ю.���\�]z�ڄP1���B0�	!����e��p�)�=a�ӐG���L?��Y06�#Ux%��uϢ���7ś�D��d�ݠQ6I1��&�H�����Y�)׫1קV$�����P����6w�������*�ψ0(�#��&`�� ��+sf�f�rD��D��+�o��]��G��t�UX{�:[�Q_���'��n঺�K�L���!�d`��}�({H���hU>�$S�q��	X�B��+c�{��!C+�@.�x]�}2��sv2�'S����	����A+ؘ�x��~cc��A^&R�Eg~j�vN�ɬ��IU��o�G���>={�!�s�A��Wot �`��\C�C3�$ޕ�<v10wbrO,���]l�[�I;fxh0-�sk���g��Z�N�tSP����}�;��B�jjCق��ն!�I_X"�L�9r�fS����B>Y��=ݛ�Y�WF����Z͖�O�6������)�\8����1��ᅘx�\bd!5�B䗽���T��:��9,�LT�����K�j�g=τ��'t��#�@�ͦP?��֫�c�cL�5����0ot�,��{ ˷�	�O�S����%"<�/.e6�~�ÖSɓv�߯��Ka)#bV�/q ��Vhe�y�W뵋6b�p�� :�$�\(�-�����g�	:�%c��,>��ۈ�D"�P�p'�8��i��b�>�k��.���FvT.Ra"]9��8=�^1h:�W�Ң<� HL���r
rGy��t�����s���o�<_!q8���a�*���������*�뒭�zC �X�- o�N�n���;���?��?�)���@�z�/�~�U�O��4JB�9٪_ϫ��ҍ�x+g�JY�ic�3��&?���Ƈ�iC������>�2;G���,����0�7"C�PU+F% �ӧH�.��Ǧ]�#Yz��q��q�.r���d���ַ1�����	��$�ҘR�yT��n6c��c������Y^�]���E~y���4b=��Y��ڬ�B��
~N��UJ~�l���U��pv���-�{0��]�o����W. ��hS���;�Dr]�H���H�_�eF6�֕�*ĝyf�ZpD���HB_�`i2�5�4S���d@s�ov[-����#���#�ұ�ǣ�+N�>*����Wz��
����[���o�%�U?t�ѯLdR���(<� lt�6��J&�����頟��/��Z�1I|���U�q��FB*���9�=�W�,�h�D5�������z�IkѴ�k7-��������o�M_�RhE_ �$�x�Կ5+�Vo��h˛��z�r i%����I��j��W��p��Ĺ�� �s�#��^ZKrH��N��4]�!#����6��>��+r�O�����5� �;Tu@ȫ���}�Q�J$�U�_7�6��w���p�gQq0�>=�E����V���=$��#t6)`[��,`FWX)D� (�4���*l~g�^��[�]�2|;�'��% �Qd�2Hɂ*�����?a�c�De�d���C�L�(W+�2v\��0P��ͳ~~�8��)�&_V�c�#+F.�
z3lT�":�GH��MC���\���� ����������m�:��+�N�x�����}�5�A�}A[�I3?Hp ��k@B�+�!n!ID��*��~���DV�g2ĜD:��j ����#�ƀ�]�<��HzJA���)v�=��s��9Ğ��Ǧ���$�x� Ew2"�M��(C*X�,��t)�ξP2C<T��B��sv�nQ�$��X��29�'NSҵ�$�3����o�&N�l�� �C������&�M��gM^z��kv)Ј�ej���
���I���:,
�x����_�	{s|�ymA�^k:��6ӝz����e{�w�m4¯.G�]|�T���k9�k�� {B'�����o�����Iv=GLo�v�e�ݛ..�>����uIXn�d�����C�3-��RL@c1+*�}f�Tr'c��ﺠ?5��"���:�_��x^\(����'���1[P�m	yK=�k��i`"0 ���J��P�����0��ߞ��+5�$�?��	��>d�<@���&�Y>��3wR�e��v*�) ��Ȣ��TŐ����%G�����I{x��I0���(8I:�JL�1��0�(d��Vnu�����#��I^R�(_��dF�r�b�07�����U�Q��ƽ�.���oŏE�N�K�c�����W��NDl�$OL䓋<~��Ϩ��i�O�n� C���۽}e�h�r�����z6�n)�	��0��y��"b��8��s����� ����VR@��`��tQ���rT45D�=^����|��E�n<�cÔ�/4���Z�OF��<������#����4]�p��=�bd�o^��,BOW~/�k�I���\Dw0��V[ù �@Z��C?rT߰U����n�8�o]�2.��f�N����ˍK�T⠓�MiBP1u	f�"�&�
O�����8�����=	v=uaPQ��/+�@�a���l�D-k�1�Wp�-���&��@H���+~\�܍ak������8:����
4����T�.�9]uv}�-���/ %�x��X��Q1���D0s8P6 Cjڨd}Y$�Sz*ol��?к!�a4�55��*��K���9 "j���":�Uc1q42�\�M!Πmvqi�!?��R*2J�Ry""�R��r]�>d��h�ֱ�J�?|Z�[z@`����n��ظ�F@�٥��浼��ǖ�"E�K_��(��`�
���S��o�JJ�`�[��视~w�bS!j߆���_@�A��Ɏ̉@w�rB��k��c~0��T�
ɋ;7�$�+*ٴ8��$@�8���K�� �j�yXz�L���|m����G�f�����i*'$��D�H��46�axw��߳������m(%���$V��⍦F̗��F�&���G�QU�c��
�Owʞ�C����ބ��a;����$~3�	�%ec��z��CE��L�$n/M�-	:�&3��%3�J	{�P�n���t�]����Aeb=��|�q}۲&�<,*G�F,��~%r+��.�"��=���4�f:p���ř`"�6��)̡Z�e��p{�m���矲q��Kg�VpهB5��^G-SaT��˅�O0��3Q��ۍu=���g��$����;�l�Ԁ�D�2���R�x	����bu#d�f��p���L��?E��7]�R~�PG\�<�h����8a`�8p����5���ɻ�WҀ�D�0 4e�h&�������ت�9(������i`����x^	.1փY����E}a䔽��K��bժ0����q�M=��V����"0��W0�s�T���e��1/�iE�s_�F.��I(D��xI����Jw�'���71m�$�-�Iv0E�����U��(G��f]���Z:O����,#M
�pW%�ꍹ�-.���b�"��X�%��}8,�OL�X�nb2P�FQ�I�	ogI�B�<�@�ڣ�:�vp�����^$R�uڍEdػ�:fx9u�s��~�xN�V́H`"��%�?gp����ϴ�Q�y���_��b�H�����=y�Ƶ���?I�x�������9�Y̧ȷIX|^�Wy#�E42|�$���u����e-c5V�˅��T��fވS��F�<������'���hp�e��@����l�͠�����W�[k�z���F�ѳuW�K���h:îن�R1/׵���Q�ߍp�`����#��$���A��5T%����
;GO�uM1��!_��>���i^�������s�dh.���M��^I�5G�%�#zMt���M�񸤂�lp��(�n�I� ����3���r���T/4��=�0�ըj����SH��Ivե_<D���oa���ÿ���N��
�o [���P���
��R����x*�HBX�)d�tQ,�	��򽛲o��k�ǟY����g������(�0;ѡ��`�i��
a���Np?�0v�f��-��XxG��ث��T��A��2h�;����K>����=z�bP��zhMj���{�	��/_e�%�I �$�8��[��)��Z�m�a��g]K2�:��i�3�Ƃ��@�\�LG�.0d$��l��G�圖�#f����@�@�� �18�Z�"�4��zVnkҩ��A�@��HG�(5��O�F���S���jS��8�mCՇ����~M:u:���Nx��;���%�8��wyȧ�!;���R����m�$#k&��-G4�7#�ˑ�rk���c%��e�1��cqm	��_���T'c`o��yJ�+��~�nΊ��%�S��k�5гӥ�o�EA�V	Jՙ�['�?a�V�u��x�a�
����� !��f/�|݋�zm�?��$9���偢P$/0evR�T���A8(.�$�RCC�xiD�j�3����;��q�f��r��<�6��/����[~�p;G�s�k�^�J��H���^�DF�6�9&����w�a���"^u�B�~)�g$A%)�=�f�w�������#�7�	�5΁:�I��8=~#(�,�ݸ&�������?�0�(A��������1�
`!�wXQ���R�7Dg�ӿ֗���W�T};C.���rAY��C:;�2�w9��=�Z{.�B}�4�~�nC���B>�5Mv2�����-Fd'�@���G��!+�	�{h?=FI�g0���&���nUnR��#�����p��1fp�~���*�ă��j�zk$��� ��$$��ϋ��)�U��r�p�����gk�v�@�'q�G��ذ� $�j�|C����	�����<a5�lA�J(��"5���ؘ���H���y���eL���`�k���ϸ}'�J���Q��D%�&ڂ�8"5�vX��G<��_{�Y�I�q���Qтm��b�A�ggX�e��ӟ�P��coBV����t��w	���EK3"�I��,H�s����;�6��8hf�������Zڒ�6 ��WS �ClZ�B�`H�����pR���}��7��%��/zB��~�Ʌ�r����}��WTs �U����c�O`ۆ�9&0 �]f�`Xk7��Ἄ�����*Y�;;il��^��Z4�#t_�>������eC����?I�	�x�<+�M*�?w� (r�����\��W]�47�� �M�y0���>T0H�y0�l�0���G���TE�5Tb���(~<]	{$֣�Tt Z)~������i�Т�C�zs�qE�q�J� ZJ��_4Y�����U�#��
F�<�����V��fOx*��f";�Y�wNWc �IY���dV	�F�l�.^���F�x�Ze%�|�a�i��\�X��a$d(�b�3�$<��a�#n�>K=��2H�P�4,I�{�&Â�?��Ҝ�eӋ�mͬ2�yc�_8���A��`#ob\x»�ş/���1�<�؊^b��쿭���%��?�By��u&�7 ,���%�?/�z#�s�_�T�s���}C���y|�n�-9 HŠ�������Ӑ��A.��]뺈
�s��v�2�����bm��
�1�e̖��&�>;�Mg�w�Lv�/���]��;.DJK��pQ���{������G'�\����sR�H�Шn޲���(Ψ��/��ÄQE���Mz9\�����M�*�#���-E�~]���3���s����
�ڳs��M��/�@��Ya><+�=�^��o���P`dtt�پ�}�9�;wu���v��tJF� '��d%J%ݲ&sS�9Z�B�[sw�> V	�v3jx���r��/�!4�!�4�~%��+��l>TC����K��aJ�:��</��a�Ε"�w*�A 㒧O�ޙz���hh��]0i�~�������Rd��.9`��rv�Nߤǁ���x �%��@��ޗ�	Nq3w"b�����#d�k�x�|l$�X@cO���iuH��ޅ�+?�G蚨���[|�=ᚻ�9����I��[��[��wy�/��_{���x�s۔���},U���gh���c���Jb%FB��9��T�����l�ɔ<�	OU��3$��В��#��A����"�&�2��GDjv�o��?�D'_������o+��qs;UEϲ(PǚR�̲�mo�b1�mz��"�ށ�Ռ?���(M�1A2�Mx�P�hi�U��MN��x�v�v�z~�V([�,V��l{�D���3D�C'oc�>�SB&g0��]��s���K�.ߢ����Q�U.�b��M�f;B�4���bD�tl�c�����o���F06._YK�6!p���hʼj�-0���=� �I#S�WR��0�Z��e�B�'�`F>��y��1�>ȴK�T (5<��{�.�[�L�a�1hl8��.�^�$�m+y��ѳ<`�l�٥�娐&ʖ����N����c�����K+��8��%�o��P���6O�?�T���YiV�D�4���uRI������Wfb�d�I�OhSX���+-�42��LK$�,K�kt�|�/�d����7����*�w�M�
̧>�@ i��n��q��g�w@(��1x�+?��;�^��/�ĢF�U�43��0��0��	�	m+�L�ObC��5�\���SY!�۹M���뒴u1<���l��E�h+��D�ai�����[�,��^�� ~=>0K$�	�T�A��=���@f� ������*�2�wE�@$2k8h�X�Y l_�q�8��R��wܑ!(��PT܀�݊
8��lX���Snv�g�1��>�Ǯh�oD����b�;c|h����2��a�%��ϋy޽����W���ږ�W�������l���R�JW�]T����o��<��l���l䃩�`�)8�-�j�	n�)<��cW"�x���%Ǝ¿����QZb���MJ�ƀ��Mp+�������|�x)�����ό�h�@��(!j�< ǻ�������m�\Z���h�¦���`�
y\@��M4�����������倗-ʋ+��Ґ�9�P~��d�˱��#�63\�`�������}q�][���`6��(�kk�s@������
��*�8�0U��/���,�-�yESv�5a!���1?�î\��*�{�P);�y��I�Eﵹ!]b����F3a��ς�܌`z����MD�٢��5�_����p*,�u��?�+�6aA�^Qn���K�=��~`.�X���(Im���BdN|��j��.�����A�?$I!�W�LU���/�4_�ҌC��&��K�ns?�݊"�D��O���|��Q%6� �������ɿ��ڝ�,�C��T�hV.{��.��ݭ�-i�V2F������-���ħ�/褜V��������ޥ>��~��x���0]�}H�G	?Za�Ř��П�r���D��9����C����zq���m6ꨲ+ثh{[�]şgC&-���/|7��/W�XE�^j�"B�tXc��4���,ӊ^u&$���ltmפ�o9w�.T���(��9t$C�l��A^�����HA<���N����%t�SP�iU��f~ <�sz������Zj4Պ�!c�R�c��5�7�2"<#Q�~��_~;�a��_=����OW���\к�݌5U���� ֱ�����s<ʭ�K���r*�MX������j8|�Ŭr���D������V���=p�U�V���W�b'Ig����,�\A���c�x��_�@Yk���#XP+��T����˜m�	�綞e�m;5��9��C���7m�XF�����LJ4���z��md#�!�gb)��Eug���sc�V���N��L�yB�	v�q���w��$w1���N�Mq{klҭS�vY�z{��p/�K�ۈ�~�T[��08!�����̌`�U&z���:�6y"v��{}�.i����>]]�ňG��d�C���o��6sɦ����!�������N������K���(IM���;���� �R.���nC��+�P����6�	�6�^4����PA@�����b,;.�����Y��9ݲ�~�)��ィ���*<��&�j���%�Z�z�r�*�zMrө"�O�v�I߲�*@���JRF��n�p�3Nh�J��]&X�A=��@�I;���S�b���_����p��~@�/-��i�v��}.f����+^�Kҗ�iV�ի�̎��=h�1���_acڻ`�#&��y�n!��(����� ��XRܿb��}4d��ҋ�2]�=���z8JV�NX&��y�k�8ȅ�7���/���DG⋮���Z���O�hP�-y�D���ml��[Q�hU��Gt�%a����$
�J�n��fw�,N-?Ѷ�� b����G�����pi�yxO�J F��|`��0��.P�Nb���p�Q{���7���R�s���0F\-y��%�I����r;���ʊT$/�SW���[��,@�4�:_^���I���b�Y�f[���@��O��.F���~�u��:vꏂM�P�.�OAF6�TP��]�` ���*E��ޢf����!9�T�o�?BU��F{��8�>�)2����ԅ������MY�`4��輰�|<s��qU��޷�?�_e���wr�|?�4s S�њI����������>�>�ld��"TV�5_Z��qz�R�bewx���C�]��#,/\��7�_�W�@���S^ѯop�]�����c��	ad˞`@KOsN��m����2����A<�u�FibL@�j4b�qu�\ٙ�ߵj��&��Ӽ/�(~S�~���X�������{U�<��H%Dr�W/-�芇c��ɜ����}n�V�mV�c��1��N����[��jXX,+{ .N�dQ����Z�f�a�0ѐ�W����2W�4
5$������n[��Qk�
ӡDO�c�;�6���2��6k��P+]��_8��+�ݲ.�ϝ{ƚ˭�K��5�CQ�5Ec�1�^�7f%��N�&t�ah��B!�RQX�w���%�K#������ �}�E���i 5�G���{A��Q����H��G�<l��X0C����a�ڿ$ᆗ2�d��9=w�N��dcaH��ωu1�HA�K#�ź땙5Kݡʬښ/��f��Y�Ǥ����_�h��#ᨲ;�LF��ab�m�k���ScXa
 Ydf�������az(/�V&\�/%e�z{�K��]��QR�ۗ��lm�b��ޕ���%���ǒ��� �`Y@�B�pM��o�ݾ��~�\={	�oGn��������Kw%�"d�T��:���Y��J��3Я������v�	����oCw7��G�Ɓ���~�-���.�V���轫�,��n��C�f�ڭ^����$ޒΥ�s��eɝ+�jh�5)�z������u��2P�Y�V��?gZ�J� ��^�S\��uW�m��s*����Y~�YM�α]_�=��c��v��@�4�]|a�B���%] F�0��A&������C��/�/�ë�0����ܦa�:y��*Ž����rf�gg��>/En��O�a�i*�����ڟ��9Q@p��Qq�q�Et���.A����Uf����0&� S�Z�Ms|rq��[�:i�8�M� �ՉI��m��l������"J��ݥ��{�Qߵ��-�?Y`��mC[C�A|��#hku���H�"$ �$թ~p�/^��Ws��'�U+�P@4���ٷV^*���ґ�ݣeH;'�b�JbSR��v3̻o����h�N�ЀD3Foշ��ݬ��p*��㰵 ���WG@�>����l�P��&۲-V������Ig���<{�q����[�����X���r����1<kH� ��Z�5��ԯ �7��㰱wTf�7�𰼽�Pޚ+|&�ch����6����pmr/u-ՂQFW*�9��P�n�XhƺC�g�ޟ�so�â����vG��p�m��O���	��QP�]S�N$��nEwX@S�z��'��Lިp
B2��?)�����$��Z�%�OJ\��s�T�o���X�;.��@��4�<U�kR�R*Q��׸��n�wv4�:+	#��O��c��_�4�UC9ܘ��7 ظ�B/v|�ծ��2���S�����r&�>[����$.�=?���1k���<��%�T�K�Z\�qW(�MC�d�ZU1����!�w6�8�@簠��l}��X���lT̸��Q#܋�t#��D
k/��ޚ���T���{6O�d��ĖKs��=FmD�` �7��5>7�C����1�-�pB��ϓ=m�_t�`-u;�ݭMzH���{��:	�`�l�`�%ړ�"U{Q�S�'Ig�����E�8A�z~�80��09�;Wղ�|U��Yς�c����
a_�M���@�3[T
�����j�鱦�(׏@�P6�y�����er����k0��(����|��ҙ�p�ܶO�_}�>��֘k�8zr�[��j b��'=���(L��{����T�ð�;���Ur �ǎ?�8���2*�)N-�ւ\�z{�u7�>"��:���2�F�
��;M7(�lfWw���/X������Ǟ.��$��~3с�����B�4w�³�Vk�?ֿ��+%��?�c�3�� 2��A�V�(����/�.�5 ����1^��8�����%рuJ<�hf����C�"�/)y����G�B[x}׵s:Ȯֹ�UW7��ǬAjFY��n�Ih(E�g��Y�j�_�.t=�A(@!�S"g��qyxLi{,g���n>բ���Z�1wr��A	�IW�$�ʞ��OC���!���va�7�#f���eU��D[o(�h�K;LE�=(�;�W
SEyh(a�!轠�D�]E��f�Ĺ#�OKӹR���9轑�h	SB=��uj`ov��dRn�F�N|�ԟ���q�`q������:�/ҿ����8@_�k:n5WsH�_"�0�K���f��0� �$��IC�>v���2�RxI%t���>`��#E�A� �� �d����H,�����8	�i佋��4��}���T���5D7X�AM��,Uo�-��J@���H	�����?%̭�L�Y��!�t�cN�����!�"�"F��^���
��C_ K���4�u����	���6u٬�ڮϜд/s �e\����dg�*�a��o5 s3�!�U�1~�������V^a�(���x�ȩ��F4�]���=��W����z��CDg����8V|�Y�tx�]2��v���t�\�	%)�r�R�-ޙ�[^�3#�Eݨ��#��`��خ�HVJ�*�(~�p~�L�_��%p�{��ö�\?���� �`L���C:4j3Xm�j˔iS\/����xF����A��>&`��i�p�� �E��/o:��Y Cr�I�;��� �)��к��2�Xv�b7_���&����"1�O��K�.���l^�te�>�35EM�bߥu^�w�v`%�x�*�Y���e�;C�j{������3�jy�&��)�o�V���ptb�(�"sg5ի#�}ѧ1��3U�UH���.e!l^4Ꜥ0�rMWJ��!�?A�žt�eF�*(űBn�E��Jb��j�}.����h�
.8'��Ɓ(I[����8fUv�U�v�} o�FL#B�g>\g;=C?��-��ڝa��_�}W��z�2%�R/��SZ)\�!I3D�fZO���o��,��m݅��$6&�����l��������u�i�v�ޗ-822��J�ϓ9i ݠ���j~&�,V�r
