��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0��sa^s����Hw�9�Y�:�E�#�BG��!��b*��e��J�s�w3�t4-�bH�T).s��B�}�C���п��4� P h�g�� ��p�3�o��?)6>����<�Ű8����@[�¶�'������k�h\J�����!g��]�h>LG�\l�
�P��x]����^j$����.�<�����=��Y��8�����#ԁ�j�4>�յ��/���B�M"�2�M&���	��Gְ�N�ٳ���ſ�)��z�A�X����Q� �[�~t�qe2��E��[Li���3-�>|L�}���G!`#���?3�ĥU�ۧ"ɑ:y_��J䔎dA��խI�i6G ����s������J���u(R=C�V�B��<Llc�p�X͂?rH����(Wn���|+�zz_ra��kInر	(b�R��em+��_61a� |\/n��`�6�k%��s����m1��+��Ѡ�Wߟ��N}҈�2[��w�h��	ר����vx��-G�)����=��<�\���J�}H�.0�i�Փ�m+>)�T*�em
�%�kw�}��z"�����R���d�Pe�4c����:w�Z�!J�Q�n���ċ�������p�ρѠ��` �7����F�6�������{�n����;���߀�Ӟ^r;6Ȧ� �cio��������I�|�;
�5
Ul;���!̟T��͖q�'Y׀D
g3��PcTJx���G���%�ץ���}F�u�I��ْ��a6��&M�N����Y�V��T�K�=T-�Y��5B�s�%�~#�\�'Ͷ!��/0��l7�HRbZ�.o9���fA�{�T����}˲�����7��C)(R�h�AC.�E�B��{#��V$-˛�����8�:���;1����r�c�#S!+
o�kwu�#&�N�0����m���"���dS�kJ1?��<�-(�� {xpÊ�]�5�,����h(�% h$"�'0�p�'֘�������.O�B��k�����F�Rzh�\��V�̀��tQ����t�$(U�aE$�}���tk��ÊK_��HN��Mi�dj��[�&ss�A����v���0l9��Y�\��C M��~f��S!ٚ��P�LY"0ude�DU呹9�}����n/����c��2��0�e�1H���n�&t?����R��V沤vx���{Q�P���EQb���$�GE����:�����L>l���۪���Os6�?R��P��2�U�{�6l��Vh�c\�l^a�������!ZS`�-��QJ�T�e����҅o���Y��>c4sU��E:�m��Z��$� ħ��)�er��sz��k�i���p��2�v�佯�� ~V�%
��L3h���	�*-&��-���t%����1x���h�!s2�;z����9��E{l?�~��R.Q���z�\�ȣ���-;��X�?C�!z�`�Ξ��O_�N>�:}e�˹jk R���Ӿ훀��ׅ9�Qɢ�8\BV+���+�dpq�c7rg�&�Å#�
�!^��� mL��o�f�A�" �`���D5��Ѡ��zC�7�z��eP��������FbWH���M4'�U���L�F��u��-vA�<�8�v�^����������i�Y��(�i|#�uYo�{:p��FT�T H;��g����pp/�n�Kz|�����|!W4T��\�w�_'L�*?����?�F��|��2�r$�����4[J;!F����o3��Q����D���c��Xa{8�A���;}�����~%U+BX"��YTP{��]��Y��>�2U�=��0a�0L�%[/��,��g0_���3ɒ�����J������\Ge���X3�V۵'����r]v=�.��c%NV��6�g3�cZ͐z_"�D���Ա\ӝLpھ�N�^ ��ny"x��g	YP.��K	d�4��y�B�~"h��r4�l�r���X����g�6��
_��l�
'���w����;���O��mN;��%]-%��,���tM�#��߰' 1/�)75�Np��"�:L��jL����ȣ��לMĚ��sR4Q���V�\qz4�{.���-���	߀o��e����K�P�{4?S�+��*z�ǾرUc���a��I�y6JF7�]h�Pc��آE�Fu�= �����N<�ı�`�P���ۍ���c�Ou��N�bh08���K�e-DpdC����c�X����zD�1�3�ɕ��R�����[��o���	Җ ()�&-�2��{�C���"�o!b�sǕY�y�qׯ������s��16h7�'��-NIn�O�j�?�&5f�\�X+I;{��U�c~�֟�?��,�T�eɝ;����ӒƩ������K���̤�3_����~�&ɝ�q�y)��=φiϣ�l+�T��N�`B�U��GD��p5��o�~e|��[�-�ai�@�p]��=������&��-Q��D���4E1'���Y���tN��A���?��;�TjZV<�CB���S��;|]�lQ�y�➘�nwq7l���!�n�U���l�EQ��T� �2��]B�^j&�Tzia�E]4XWg�YTm�G��!���3�v��7;�!�������LC��� ���?��e���u�x5 V�b� H�Ink��|��-�7����'T:vIz�88~Z���o��X��0�ʋ�ũ�� �F�÷u~��G�V�r�<T�D�@�d韁_<�|$�Em� o�%,�m��)9�j��ȷ��TY�+!�S;�15�_�9MO�a�>hS*_vr�R[���Ec�\�#P2@*>���囬KZ>�Y�=w�p�y �������ݪ��!䩾y)�V<��h*>�bI��?k���N�"~&Ib	�n��c�"�@�16����A0y�=�h�_���i\��0�@w%s���@�/�5��Zn�şF�ù�7�+H��J�C��'a�H�fC��nE<�(�L����]=���[��:���ƫ��/� l��V#ii1����B��*�j[0F4Y�����ԭ\�������X0�J�iJ�ϯ��׀�2x�b�s\�������ְ�|=(��R�O`N�x�����Q�L�1�fgs�<!#�J�#�ު@�Аu�%ZS[�#����Cq��Ź�8އN�A�)��>�6��x]Ҡ2���[�M��Si���Y!*�s�������O9���	ϕX�m�<eƐ��XÚ����Af׆%Mp���]K�����  �g�/�������g�ݒt��ȿم�݂��h 2����b����^�i	&`���`��9�5����L�J����/��V �q��
/�HEV~�����;�r�{C�̟���<�Qy§�(w>���ZӺ�@�ls?�a2�3^��M��ú9��&�K)e�w��]�\����V�Y��t�R����ύ��5�29mg�C�����������=���eg��1��P/ArQe8�17�N[09��)X��҇�ڣ�Ў����w�g�v���j+�t˶�ϝG�7L�n(7p_��w2�l˗��/BM:<$�Ֆ�B(@
�)g�t%G�*h'ɤ	�������o\��oP���#��L9�J��U���ϟ��DK�s�2h���߉���7u����~$����p�w&�3W$ݖ�ş�Yݏ����kX.��"�!k�Q;�0ѱh��,��GW��>�9C�S���Qůׇ�kVLםN���b��Ivv�e����`i��[&hgo@�n���kq�\	̯�)P�*���(��W$�U^�fBL��1��w��	�s��[y�9y�~��]�A��}��$J����U3+�(وz�6�4�J/�W�e��,�s-׿;�A!iC�ח��▮�0^����Z�� H�2]��\��-JW<~�����y{�}@��=~��,�D����kC&������nd� [��3C�l�_�bkN� �)8O̽Iw7.�>ǁ�i^�c�3Z_���1M�&�<\�H=��w���6Ö���.��;O(7�^�^��r`�d���f�=G���k�bV�o'0�T��]ofb�{�<7���_����W��}��Lp�٣{��f��5�儗x9��ٕ�g��ft����G�@�f�,p�G�>�������!ڡm����Y��[�/�y���r]w�l����HK��p�o�L��G2���b����#7+s����$oO=Ѣ��B~��������P[-Rv�g��d"|ǃ�ự^9<r/6%��>��� ��*:�ߧ�u��C��o�3VJn$5Q�|.�&Ȓ�ỷ��rC.&ӉE����&���+��Ъ���z�[vt	�'��)�/P�]�"񿵙z�1���x�h �L�2 l(���7���d�|�.��C�m�~(�E�]0��VI˖.��2���`�";��l ����m=ky�6�s���W�Ut��0X����3/@�Iz�U�XO�����>�d~�?ooR��k�Ani�C)W��/v�<���:����Kn#R�A����v���&��j��	���{H��z��x��]��,p7��k��?;L�Y��ҵ.$�%�;����H������S�J9"��f�	��F�q�?���>2x�K!+��H�\J��o��nC��#�h�+�G8�EN� ���ʪ�;���?ZH-����V���g4�B�p0�&�M�ey}au2��r�a�<p@��qyw��Qt���29/�$E��O�w;�پ8�Мs�V�jv'�<�E+4�t���d���v�A�^_Q��;b%OV=����'��P��G�g�/�g*o{��ι����
�N����	�@ι�݄����\���/$B�z�ꁿ��5�X��ʿ�z)�M��Oa9���h(Db�:��6��洑y.=嶺��
��4k����}6=�p@�BG�W�G�w��|i��2sC@�İ'!��Ǵ���n!��sn?(���4��Q���{%�d��''*= �7x��V�ݎ�EgO��[�7��Jݸ�X���x��uj�u�;�;ނ��ޏ:<�ut,���EW;����I�#Cޣ$�k=�,�:�5�+�[m����++����Q���u6��R}�
:&+�}���x����LXw��T������k��]�R_�_*%Z������p�f�t���Ǐ���}SKv.tKS�@{�x����9��f�>�n°0�Q�:�B�׶����4>?Y$	��vM����,��L�h�#N ��g�~)�Z�& }|SkZ����y۝��P�1����1,��g�w�>zo��Z��ۛ�>���?)���,����A���[�Џ�C���\�yĥ���:�����.�(�9�.0�����*����<K�Sn�@�?�����xs�ù �&��bbw�����lS���(Q�ݸᇉ$)��>���R� ?à��Rk�#�hسvfJ]A]`�)��$�Ӄ��^a]U��l"Z�W��.�L#}�J�b�A��D;t��MDJ��O�'}6�F�$�`������ˎ����c��Xj]�%�zg�=�B�Ip�
�F;S/��pp��d�IJ�꫐	���hǵO�&nO�T���� �`�5�y_`Ї�L,�5�ؓ��"�}����4�6�[�ˋ����6�J�Y*#LEO��Jv2��T�0�8S������~a�[�ň���ޟm��)m~��Y��s�c� ��}v�����U���:�n褤42i�/��G�w�%�|��WoQ�f�:�_�`�G�RC��]�Mõ܆z��]�,��.��3��d�d����t(�l�Y�à���v����4�QM!��
p�1Ϛ�#?0�}��@CY��H��Em#�iç]�ms?D͑����:�y��zֻ�����B���GD�ʂ��������J���;��:�d"�[�X�C� U��S��hA�D�	�GI�e��o�mE䇛"羥����~.
�˱>UL)��$w`]�qփ3�i��n�_Z��D� �W��W8��{*tg�uC}��%��꺇���.�f�=���dB�zUL��� N�q{�d�9��H)_0���GE�F�;	��Z�ˬ��.6�P�6��uF�g�����z�ܴT�F�;?�z��# 6�G�c�xQ��/I�^�>h������*$$'�l�LTqf�@��������)D��rWu~�ͧy��	!E�0ï�Sa�'�p�Q�J�ρ.����� �2�+Pi����+����w!L��X=����p+n"�(h�Y���H�$G�js/����bA��&]x��l�p��F��?Z�!�,H7���a�Q"����J�,��Zs+*��\�,r���Ipڀ�f�eߩw�7�j@�����Dz�H
ɔK��ԺN[�шV/�s���
b���LO�^u���2ξ+}���W�SE��I瘘�,�����VW��]�k(	�)���G^򾌯h�v�H}f���_P�0y -��/0L�	^)Wk�
�]}uB��$�Ğ��B�����M�f���.��>�dk�osC�V�eQ�Wj��Uh_��7rMW3�6S���Z�w���#GL�G�<�bށL���@�`�?��0{̀�T����3�{�����TcQM[|\����e݋p}�A��4��/8�H�b[�����.�����i\N��M�5Yu����-�2�Jnyx�О��M�?�c�H���''��r�E�T�=J%�O�<l ��@����<F�����Z��3��98(��^���y�M�wv�H,�����e��	p�v�� �y@D&-I���~��bu	�9�\��T�����`��@j�͗������s����Ba��&}�4��Mn�ˀ�avo���}n�m���/�e�bYvU��V��d���*]B&Ӓ_l�"����(R�-��"��% fǀM��X)�X���,ۋN}�*����Ra��%"��~�8��(��#��nxbR��X~�-t4��u!��I���$�o}��D`�����-M�T]y�O��ݗ��D
s��4�GO��{d"9��x3R���*�Qsåߪ��d�vhM������9ҽ0fZO�U��i��,V�e���Fѷ�O{�dph��p���|<����0A#�#j<��𚤗th�����N�p�Ȥ(�Pta۱4Ş����R�6KϬ�Lj鮁 a+�Eڬ[��ߕ���wR�X{�7���'So�����A��NU���u�����.A��Ҕ�Oϱ����(+5�0�}��������N?���h�?=uc�e��9$���NH$�+;��ܯ�̐ۇ����x�����-7t�Pnv�U�X��X�,�kTY�Ȃ���}1�u�O�׫)y��V����L>���w8M���-�y� 9p'�U"X��?s��~�\�e�&�)��c~hw�8;0���7�:x.T�[��pW�{���2qarKB"ie��@?�'+���f
A٬f[��$+����*Z[��v�q(d�^�K s6�f�W�e=�c��-�>���ߌwV�K��[�������Zas�W[.�v�*�D���ht�ee䑰_�fDmM~`���b����8��B�� U�ǩ�KGO8Ò�+&� -5E&�d���Q�Ύ[�$�j�f�L;W��E�����uf���AG�|Sz@��j �ߙU,B04�T�}�_���3�4N�U%�������1�\VA����inG{-���F����$�	ࠛ��sg%� hc��:Qi�;�Y��j��Z`���F�7�0x�ׇ��۠t��-�Yf���K����Q3eK�QJ���'��k�2Ѐa�������5G�]�KxIVδb���C�#�����{[!�-�v�Y�MT:�4R
�7�@3�`> bi��۽�[#�a��T."�
���xG���"�O暈�CL�׷��'�fLĈ}k��rI qqڒa���O���2��4'��A,�/���1:SD&E�}��̊%���c٘��CaOQ��E�}�xCN���?��6lI�F�� HҷӸ��*��t���'+)�c
�iV��0��Ƅ�_�a��a6��VA[LZR��-{+m����[ =[�@/2g����Dq)Y&!��(�)��i����w�gaY`�y\��MB�zG;JTBA�~���
_P��DJ�o�`�@�?#A۵	�^N�ob�h�{&����(@�i]��鿍=����q�<|ˍ&�:ʚ��(ߚ��}m=O�,I��.1����XL�������34*����ģ�����ʑvY�?�0��j(v�c������D�q�Le: �yu�3�*+�D���m��x�ڲk�*\`��,-�FAĖ��,�4�H�zw4����WF�����=''��E�<����|j��|�MeW���&�[)L���:T�\��Y���
I����q�B���ѽl.�;<�8m��i��U������j�'�a�,�YcÓD�R�I��V�B���M7�����^�P�{�d
���aq ���<\6����ӑ���6�7s ���\��U6��P���t1�s �r������,w�/mrfݽ�*�lv!8�)䆵�5(G�RG�u졀�U� �Ueq���A[4�e36�;hδ��B��i���%9''XZ�^�`?`7�3g�)�b�ޭ�����s��%~��3�yM�`�������fz'�Xu�cFYM��qCڂ:a�-03ɵ����,V'��o��֬�j)�C�c�4�|�1Υ���A�-�F?ap��~T�+x��-{�=��b��o3�s� .�
Z���1�b ���5^حM�Wi���ei�g��Bf�{��3 m��Q�@�/�u����,�/U?z��c��X�d�j�2^ ��Zs�
V�D��)Ѵ�ʞ+�k�/�c��t�ݩd���M$dx����s'1T� ɒ��Ѧ�8����y���NV�3-���{�g'���o�����^�FA�eTiDQ�[A{�?(����0!����'�b�����f1�? E�=����P���SE�mzd��Ou|�<�0o	�r"_���r�Y\�:3�s�"$zD���C�@�y�Z���$�4�}�����,y��N͞	1��+�a��}�Į�	 R5=��
��r��Lu�[�A'𹾪D0Hr�@m�C��g3��ҙ��H�J�]�F�|��~�_\h�	[�߾�˯�P�x���B4f�o�ߖ�F���<��A�O_{��0��^�^n���wA^Rm+�Qv����k�p+R�lq�A��ΉV��I*�ࠀg�d+
��ZY�x�g
q�2%o����� U�	��G�����#�����P{�&F%z�E�47,�WHe���/]�*�Dդ��>�N ��$�:/�9hn�\��(Q;^������K�b[5S�3͏���D,W�c@w�0�zc������Ae�~��"_��ߣ� 4�Mۉ�* �^>��G2�uW'e��^Ɂ>Ln�B������%܋�򞒘�) $&!J60煓M�%f�߻�-�516CI���9�����n�j��J��Ӝ��U���o�#�X���	w\֙���CD|jH�<�0MNA�Z0x!��!�(�P����\�WI��ABJ|�FY�d?��|�K�/L��2�r�J���|A��� :}tR����rӹc���U*
Xu<�]n��aH�S���:���!��ꋐ��a��=����K��?p��c�X��f�5u����	��uk+c��,@@شIm��J@�CZ�q�	��QG�lːy�E����GE/鏣sC�ء�''?����w�nF��Wۗ���+�=�����v��M{���ۉD�.d��Ю���6}{Ц����X��z�]��Y������5N3�����<�8�i�1ta����97��O&횷�b�陏-*�`	s�(&��	#���(��A���`-o�<YK�f������" �Y��+������k	ۯ�gt.����$s���c�� u>��1m^��7��5,�(�/�98��2L0��I�c�^�(🍖J0����5b����Vt�"'���U�dӮE�'�G��y�����ٔ�7�		A9~���==Co����E%1���W*�W��h�i{	��t
���a��?��.a.���N�L��<������3!�ٕ�!q��/u��y.7���vZ�"��0�� ���7�'n��^��H.��x�1���j���&��*H�����}P������Ԃ��P�"�&��b�n_�y�N�a�4W|n�
!�� Ue�}��sW9������+S6RW>�:��b�V��+�@�g�
�RZ#Bӛ�Xr��Z�����}��M�DF7�+u=�H�Zg�3A��5<��!s�]�͗
���4���J��0�%v�ܣ�X-������q�h�{���]��>�YiXR�>J��j��=�a:0�-|m�5�"��i�߃6��������*�pQipNZ��+�g�-�q�Dɑ7S.�(�E�1��ץ̞�vNq�R*��0+�!U�s}l�w5+�*�V����v�B vA�*��hY���V�ҷ����?��#Y���G�wǜ-m+i�q��|s)�0x��bO����LpF������x�f�S!�ղ�*��7��7��g�
L{��3�>�h@��\ E�d���λ��kՀ��JI��[m����`j���x(5X��cgYT��j�7��٩yt@��u���m��^U���^%�M��T�	C�|��YbC=yRPQF�׊��,�g������^�GbBs���
L
�Zr�~@�8E�'MZ�m��*�&��)D�ٖ�v�k%f<�N:�oe%PQ<����b0@7֥�>�B~7�2�)Y�	[�G;� \L�%i��3L7%�V���o�XJ�g=�/���m!���t�څO}���/E`�7�b�M����T2�����G����-9�Y��O ȑ+��wk�4��(�a�YD��W�:zI��zxpa�|<�m����3(��A�U�<�'5B���f�YJ�7��9-��ҁ�4�_QJ�t�sוB��Y�@[U��-�l\)b~�He9�jMe\f���7��S[��G��'Қ�ف�#�~Žl���~��zY���zщ��x8ػ��~�>�=Ta�)���t̵�g{��³Z��Q�n4ADQXo �ZF
z�hp�gp"��1����w�H�h�\SӅl�r���[����6�gՎ~7ȫN��2 ��֟�^`��鼊�� ���8���/���PD7֖�'`)�4���L��\�G�9�q�:���Kb�V�wC�ci"U�s�7�2>=�C/'^~Т���d�%4!5�[�ѫ+�1��(U+.�L)��X�B�E*��@qR����p��'i�G�,F	�icN�u�۵�tf��L�u2؉�$1c�g��C�31Im:�n Z�z�QA�c��*�`�0i��M�K4[��ޥ4B�*���mE�6�4��7�;�����S�tB<�
�Hئ'Gh]*s�ϓ1냛��c
4��"�d��hm@e}��cU�(z���I�]/zX�
�'������5��U)�.=��Ճ]%uԬ�[|`qB��\�{9هl
A�)�Pj��GG�p���݁�y�����8H5�Z�(o��Vṧ&ⴝ��?�ƣ��V���h��`һp�"�ņ�?V�H�����,�k5ԗ����N4J@	 g���A�ۊ8x���W�*ݝ�ir48s���m��9Ws^B��	�K.�U�=�a�߿�_��W�j���&�x,��Z�H�x
f.��`��x��R����ja��=Sn,Zv�Smm�ꆔHD)nI,�<��ZH��}��w\``�G�T<6ƪ�7E]\�--Pґ�"�v�~F��l|u��st` Y����'�kθ>y�f
���Т�RO���췤ë�ڏ*��E�H\T�P�nF��o�V%V��*.wI^7�K;�W #����� �̖y�-��!a��g�=e��"�M�qR�)�����3��́r�O��*��ܟ�s��g <e[��
>H�B�+u�<�a��\+2�a�%���>�`V0���D:��������{�<�YV�A�7K*ݴ��C�z����I$|�}xv1���~�n��t4�ow�6<[��T����*���U��a�)|>�#I�İ8��Ǒ�H���?�Y&�n��5󣘔9�uJ�D����BM�o�=�W�ϣ��f��M�iG{�&�(������tZG���yA!��H� ���o/��J�3%TCך�K�|O���f�\�
h^�=�L*�3�>OT���\8o1m�!Yn\��Dh�cD��c+��
��ZJ�*vm~$;��\��L�m1&�Pf���Ai��/V���.j_�O�	����KE���������HS�O�&�=�t%,��fꄼ�h{0A���z)~& 9ǿDZ�U��C��.�����UW��_X���.�&j�W^(xhY	H��y�I���؍�kZ�wF><I�ؙ�R�RlN��6�#Dg�?:������B�x*V��,�eY$��-z��D���T"1[�}	`��Z�z�'�.��E�ڱ��d�L �4�N�Nа�#�ۮ�`"h��S�\��0h
5=p1�KJ���a�/5y�v�}zZGV8�ׁ�<z����8TO�4F��l�oس���6�	Z^��`���0����࠯�X+`��}vZU`R
V��2U�q�UG*w孪4͕��
�Lx�٬<v�9�Ųg�Š��u�]��}#a;GV���qUi�*�>�J�D�����x	l�����SF��<.�
#�<bt~d���X<�&G���3��ju��`*v�_�Oɴ-�c�u�C�}��o�oMA��7W�J��ݱ,p�;�)6a�NPUB�5������V��q,�lg�g���1������/�����wa�t��������c#hӐ�@G67�P�\$`��;H~��x��r�g�)�k�&k���Hj��+[A���[����Y�f��k��z�KE$����lw&�b�t@؆�Qclt���E-��ɝיcB�}���q�o��qjB��FQ	��� �*aB��	� G�.] ���3��]�kI}է��ǉ4��]'qG
C]����H��cd����5���Љ,{U�r��<$����(o�9ld������P���T}�tw_������� ��/�cF$s�����On�VGR� 	�
* 	�|s :�M΅B��S��w�^�ȼ㒔�`����$)t /`v�2�c�����Q��yFЙ$����6��"
a�,(C<�Q���LG1n���r�I�*"�sRX+(��R�C��A�~����"�6� 5�3~�?+�0]��_���nsJl�Аx���yd�n�Ɓ���v�o�t�(UU�d���P6�{
�ߏB�
F���c�.��r�-@1��[�w]-v�G ��]w<A1/%��!�ն��>n��m ��Ѐx�n/迱�z� ����yID�|�O��P��V+/�gRr���E��
`�C��=��N�)'5'�r�9���7ʝ[L�hY?d��m5Y#�%eT
���f6_�j@��0�[s,�[H���\%�[�HŅ-��o�W&��5�.Bg��	")����;Pky��Ӂ��4@�����;�PF�6�>N 8��W����ȽI��lŋص�]���^���c���LKڑ�
��9�L�'����t��b�w3H\/$���\y��;�?�.�g&\��N�~P�-����L��;mc��k�ȖJ� 	���^��˔3	��i)�]�G}��zl

h�B,j���7=�z�Z\.�1�[̻&�������g�D�I��.�\7�t����>����%�Y�->�+aq��<�	4Bai<u�oun¤� �x��m���T�k���GE��{�NsĂC8����!8?:Ij���� }rs`� rrBf�UT�|�8��&v_��j��1�h�3�e40A�(��|x�˅�$(%hq��|��r�rnq,����b�Q��`̌c�����hn��3"�N0��ۤ���2K`��poȞ��=_P�����Ls��GwG۰�~�~`��<k��8a0����j�6����S�o?�e;l���� ���P	���V|���x��BC�{�N���=����Iho�1tΛ�K�Gfޙ{�3rMl��]�kt�S$H�����[A��w����)��	$u	��#tou�9���?$��ڭi���CY�G�`S��#����d{2���̩ �X�<�DuQHu��;e3\�e��R弥�a���v��)�d{�R�P?>gko���@{�"�dt��_�+P�B�t��h,>P\�g�X{���r��Q�yo������]o��Q����j���k��ڟII�����>l	q0T�0�g�=4�?p�:��+u/�.O��R\�zj�ר�:�IV8c�:9݆����Nxsܔ�I��@�����NG�D����Y���1�� E�� T鑎��VҐJ�߂uW�}Z�HU?�:
U��͖��i���;��TR�ʪ��^���_̵�s�Nl�6O�9�~"(��@��w��=�Жj+�z�b�%K��p;��L��֧#e)��otM�(�t1j�.�[�1�g��1�y��֪f3�7h� #�bD��'�E��)�P��#7��7��Y�����Qi.��yJ�c�ч��ǈ���7D����N^�#���x��?H��S�	S����Q��ݭ����+V�%��ĺ�����8����DxoGI��#�`�x�C���vq�+����
�s�vv����׎�C��~J����s�H5����Z���������l������{tX�z�[�����K��q�gP�=T<c`���!4?�;�qO�6���M,s��\.��z�J
k1N���x+�P4�HN�@篩�|;����_���{�y�WE�/�C�"��xw�i�^��~�?b�5�B1n�#�G'<���*��QD��6��L�U^2���X3\v$�n����S�����Y�񛎑����Jc��3Q���K�{Z�Ď�A
