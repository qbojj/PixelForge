��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����o�{����5�{�GW���Z>�/�'�A������ƺ%�KEL@� �I�)��d��:!�/���T\������E�Q7���"���D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����vxU�|�o�0T�!(꣢���A�Y�:�y�lPJ%	]O��˰go���w�2&��xc�)-���~yf�6V���qt�
����$����P���7y��cg{GR�Y�+O�E�v��"nTё m��E�k�~�-6� �#�[^�������X~�;b�����QFg�*����9*��-�/	Qy��o�7!��
��f_N�cN}�O��k쨝��F�'�l�M��4��������k3r�u��K���hw�/&�����Û^�	��r�E������R	�C�8Td�;�n_����J�̌)(� �``u�����]�_O����%
W��d|޺;6�̧@��EἹ�jD�)(�yn�_��^��
0�c>� ;3T`>Uf_¸}�ԝ��+|�Yo�PB�m3~n۪�b%�߱K�;����i��?��,�[���!�q<LFv	����R^�Ӝ�����_�4[C���4K/Ӫ�L�V?�yb�7(K|nL�IǑ7Q�%�:���$:�+�90�˝0(���!�̧牪4hԅO��^�2Xw<���o�i����ym�v�/H �"�4Yb��[�/�5�\���[П??�
�P/~�k�ȱ�B��]���5��;�WZ�l��R5��͞"�2Ȼ'�3�}�%G/�l�#��J�6�U�V=�J/��+wQNT�Z\�Ȫ7x���!��(���8�a�4�LOeY�?񱋧ʹK�}���d��y�D���2>���iZ��H�)���1/c�ܥ�Ս-pl�XK����n��A[7�M,��S�uB�ۆ���J�@e纟U�p�p�"�����7���I���;����iP'�ټ�u'��x8��>���
���SeZ��<��h��m��P�5O���M�dK�YG�*Qe�A�}zp�E���g<4��B`�@��6���ԑ��/�=���n��	 �:5Ź�lX*
�3u��ܫ�&�����U�d�#;l���9.��?/�ɪF�ԥ5b��k�����n�W}�`�EH�ER-j�`h��A�p�R^�Hi�B6��|s��h�`�(�92���:��ɱ��m�����ȃ&{g�N�]37
�S��s�Р}ԣ7m���qܞ�RK����y ��!7q�Ao�6��T�ü$2d��Y��ǳ~r�,��+�q4YjQ�/>~@�k.���W|��m����鍭��i��)$z���tu
�����7�D�;�2f���]�K6D.�P):���Vb���8V^��2�v5;=٢Yݬ��So������Sa��ڬ�}�_�oV��LIhq�q�A�f��0�ʑ+m������B���L
y���^����P =���dr�*2�vÓrsr���/��G�_�;�X7I���J��t���҉.���L�}d���M�_*ѥp��݆��E�\6���'fYWcLVŬo<�|�4[6z���"k��J\�.%DJ�Ymd�4����vPQ�lX����3"�c�Xl(J�C�-ugaF������S�h)ʚV��%�!Dw����`��e�_c�������f'-�Qc�=�+�o,V�U�2�������H�M������`g�	��+P�#rd����
1T	j�.�#���*�����A/J������#�ncQE��@�>�?�ʽ�����ǆ���D���3�4Y� U�l�)h��`<�o�ݸPV
��i��^52,��B�����4���뢯K��M)���#�ݷne �y�ؖvh�Y4���1�l#��-�:Z4wa� @�p�s�-�.܂H��c
�]5A���1�w)d�=�s�D�6���{�[d�2����R0i�[�k�i�첥F��$l׌F�gz��b��I�nR�;>���4}%l2�5�L�j7;	1}sҳ�"��&�<���w@I�p#�s@��]9cY�6n�f
��-���2G�]�#|��8Սɲ[aҌ�+>��@�� ;\r|	ᇗ�u[6�{CO\ꄱ��d #[LK'-ՠ����F�ܞo�������8:�Cb�>&EU�]��r��1BT������G�`�y��|@!�UO&9>X�zZ0��:Y��М�l�nؚy˷����S��ǁC.a�4/B� ���|e��vz�A>�grx�ǹ=�����������/.�$��Gڒ_�Ɉ�*x�wg��������fr���x�/�C���H����E���_=��2�_�;�:�Zm:І� |�l0[�xY�ڟ�W_~���Q���P��2�W�WH�r���tf_�9���)*%q �^H� L�Cf���4��;r,���U@/fB�a����U���e��c{|�x�]�o���:�t���1��f Q�A�a�c����L(�GѦ{.Usb'��y���ed�D������N���8Ɵ�2�Ie9�^k�ϋ��ۯ��}�<�����4�(a4o�ɐ��7)�Z��S��t!kyYwi������S��P�X�W@�)�ؗ "��fE��Հ"�3��C���Ux2��_�0%d�ǄAp`��Í�������$���b�U�֯N�F��Y�Ơ����yጣ�o��ߝ�L5���1q��u�7��(` }�`C%�t0�z�y9^�'�$�g���a�JrNI[;;�~��#'G_�[��k�$$!�$���)1��r������$W1(�m�&D
<��2: ����Yu�a�o����~����9Y��@Ճ}��D������A�
(�M ���L_�H=�-žۖ3�A3��=0T��BO��ٕ�۝�z[�Ӥ*P��*�.qtz�4��$x9��"1��;��(�CW�LֺH��/�|K���'��|8��c�����~�zx��za5d������MbW�r���0�$3P=a��Z�9��r³nh�";�{s'¹&O|�PNM:*(��U+��qv6���+c�C�6m��Ɣ�U+�j��Vvx����i�Y�S��}ؕi�Wx�B�ק�\zrK�[8r�@vI��=�_Ŭz9S�q�C��L�\/�4@��;R��)h� ���_�' �/�	��c�(l3N�w��r�Q����0��Eˡ���..} ��q�	UdB0�1]�֗��L�֗��nLĂi�x��7��=����Vnב��De�^_"S$8�~L����cȑc���P�gj)nA�P��Kc3:�nl�sZ���D�nf��"����%���=0�u *���R��������$�ķ��� A6��do'Ξ��Y�yJ0��������d�Z�ڃ���qt��p�t�X��.Ɂ2��+���9o7�8�(�3��QD��@ii;�EՇ*�Q����K�Q^�)?=��P��6��@#�`Ȯs�WnGo���(�E�k͖��J��<���;�k�E�1�5I|)�+	n�6�:�B�T.�C8R�*���w�j�ݗ��j'��}(�ec�����Ew�����d�0�~*�%i�5uH4tQ��8�P�(ƠT�-��N��뷤����%#�	R	9�s̞Ĝ��Э�n15��X6�b�=�����R�1�l��d٪�<��<"��,B#9�*�Sh�d��'(-U���kA6�&)�|+�s���$nvP���m��vQ����p�g�=}�h7J���iV��:Ŵ�J8GC���BE�R�g͸���GZ�����X=}�4�90[6�����c~ {A�E�4E����kJ���Aw�I�Ѣ�cmܷ�W����������z�d��3_K3�Z�T�*��ѥ����;���U|%b�S|��iYշ���1��$���XTY�@s�ժR�tq~5� �H!�|����w�&��M�u�F�q8/���8<���|ꐋ�S҅�f����`;$A��vx��E����R/���*w��d�1����&�`�lȀ���uMQ�<dS�e�A1e݇9,!�I���Z��������p
Z�$��v��Q�o1JZ��1H2MiR������Q�g��֐��f{�#������0���r��c�S���C�Z�9��(T-�ϔ>����7r�wDC�v3�}pZ���b;�.u��0���."��ՋA�; g9N'��V4�H�;'±G9ȗ�U�)�!=(�V��!�P�9*�G��m���|VX���-	��߾�\1g��0�֛�o�������D�,a��ۺH����=4��_�+� ��F}�p�A\��ڝN]�e7�d���b���XUSF����8W�������9��x�y�<ߎ汛�0��X�ո�CY�?gW�x��V2���]:�&"�po��5�2f��\J���%1Ȯ��7��b>���\`��z�������8kH�(��#�/�槠�/� l�eFM�.�Ѣ{ʑ�.a��	�  * �qr��Ё7VW��$�A���������'��-�}��39M��R�]�+P�b�p'EM7*�O��SK<��Ua�P��E�#Rj�L���&F�Y��/76Ae�<�.���j1��I������w��%�r;ٹk�s�0�=7��,�ǾH-���f���[[W0QZd�+���o������&F�5q�,i4�=ru�NiO  t�QQ0a*������Z1�r���C��+
�h��_yZ���#���`DHΔ53�@�����v�օ5lE��)=&��Y$X�a���9,8�)���v�-�<C�Ceb\ۋ2�jW�����6t��jI�ΉHd�M�������^$ ��?J���X�Kb?���J��=���P3Z�ʼ�Ey��8Qa�a����X�6��9/Lc�\ d���!.	����^M�P�5_I��*�l�.!���X�J�o��y��67�8�l�ZZ��fƞ�t�Ŀ$��Э��?F-ϋ�/��	+8�'�}��2���G��zRSg�)�V)��*:��t����j*@��	��~c���e�x��&IZ�c2D���bg��u�8�}kǴ��.>�1�T��&��=+���0h�~p�³�KϘs��0�C�SDt���,-�A��fm
[�`"���x�8Ka���M���G��hk�
���z�iOt��W��|�����ͯ��������Ε��:ex��gp��@f�r�Ȯ���&�2f���9�3f>�l[s���ZpxwhȨ���r��5h*+��^m��gJe�w�Gv���-�鿝w��0�1�R����ɨ�U6��S��@~W^� 5,�,B�)��%勋W/J���i���S�f��˹��:���v��ψ��֏Fc�?�$ےЊ+qֵd�
��q��0�zO�d�I�O�G���J6���
